magic
tech sky130A
timestamp 1697586785
<< nwell >>
rect -115 2845 525 4130
rect 675 2845 1315 4130
<< nmos >>
rect 5 1475 55 2675
rect 105 1475 155 2675
rect 205 1475 255 2675
rect 405 1475 455 2675
rect 745 1475 795 2675
rect 945 1475 995 2675
rect 1045 1475 1095 2675
rect 1145 1475 1195 2675
rect 5 -45 55 1155
rect 105 -45 155 1155
rect 205 -45 255 1155
rect 305 -45 355 1155
rect 405 -45 455 1155
rect 745 -45 795 1155
rect 845 -45 895 1155
rect 945 -45 995 1155
rect 1045 -45 1095 1155
rect 1145 -45 1195 1155
<< pmos >>
rect 5 2870 55 4070
rect 105 2870 155 4070
rect 205 2870 255 4070
rect 305 2870 355 4070
rect 405 2870 455 4070
rect 745 2870 795 4070
rect 845 2870 895 4070
rect 945 2870 995 4070
rect 1045 2870 1095 4070
rect 1145 2870 1195 4070
<< ndiff >>
rect -45 2660 5 2675
rect -45 1490 -35 2660
rect -10 1490 5 2660
rect -45 1475 5 1490
rect 55 2660 105 2675
rect 55 1490 70 2660
rect 90 1490 105 2660
rect 55 1475 105 1490
rect 155 2660 205 2675
rect 155 1490 170 2660
rect 190 1490 205 2660
rect 155 1475 205 1490
rect 255 2660 305 2675
rect 255 1490 270 2660
rect 290 1490 305 2660
rect 255 1475 305 1490
rect 355 2660 405 2675
rect 355 1490 370 2660
rect 390 1490 405 2660
rect 355 1475 405 1490
rect 455 2660 505 2675
rect 455 1490 470 2660
rect 490 1490 505 2660
rect 455 1475 505 1490
rect 695 2660 745 2675
rect 695 1490 710 2660
rect 730 1490 745 2660
rect 695 1475 745 1490
rect 795 2660 845 2675
rect 795 1490 810 2660
rect 830 1490 845 2660
rect 795 1475 845 1490
rect 895 2660 945 2675
rect 895 1490 910 2660
rect 930 1490 945 2660
rect 895 1475 945 1490
rect 995 2660 1045 2675
rect 995 1490 1010 2660
rect 1030 1490 1045 2660
rect 995 1475 1045 1490
rect 1095 2660 1145 2675
rect 1095 1490 1110 2660
rect 1130 1490 1145 2660
rect 1095 1475 1145 1490
rect 1195 2660 1245 2675
rect 1195 1490 1210 2660
rect 1235 1490 1245 2660
rect 1195 1475 1245 1490
rect -45 1140 5 1155
rect -45 -30 -30 1140
rect -10 -30 5 1140
rect -45 -45 5 -30
rect 55 1140 105 1155
rect 55 -30 70 1140
rect 90 -30 105 1140
rect 55 -45 105 -30
rect 155 1140 205 1155
rect 155 -30 170 1140
rect 190 -30 205 1140
rect 155 -45 205 -30
rect 255 1140 305 1155
rect 255 -30 270 1140
rect 290 -30 305 1140
rect 255 -45 305 -30
rect 355 1140 405 1155
rect 355 -30 370 1140
rect 390 -30 405 1140
rect 355 -45 405 -30
rect 455 1140 505 1155
rect 455 -30 470 1140
rect 490 -30 505 1140
rect 695 1140 745 1155
rect 455 -45 505 -30
rect 695 -30 710 1140
rect 730 -30 745 1140
rect 695 -45 745 -30
rect 795 1140 845 1155
rect 795 -30 810 1140
rect 830 -30 845 1140
rect 795 -45 845 -30
rect 895 1140 945 1155
rect 895 -30 910 1140
rect 930 -30 945 1140
rect 895 -45 945 -30
rect 995 1140 1045 1155
rect 995 -30 1010 1140
rect 1030 -30 1045 1140
rect 995 -45 1045 -30
rect 1095 1140 1145 1155
rect 1095 -30 1110 1140
rect 1130 -30 1145 1140
rect 1095 -45 1145 -30
rect 1195 1140 1245 1155
rect 1195 -30 1210 1140
rect 1230 -30 1245 1140
rect 1195 -45 1245 -30
<< pdiff >>
rect -45 4055 5 4070
rect -45 2885 -35 4055
rect -10 2885 5 4055
rect -45 2870 5 2885
rect 55 4055 105 4070
rect 55 2885 70 4055
rect 90 2885 105 4055
rect 55 2870 105 2885
rect 155 4055 205 4070
rect 155 2885 170 4055
rect 190 2885 205 4055
rect 155 2870 205 2885
rect 255 4055 305 4070
rect 255 2885 270 4055
rect 290 2885 305 4055
rect 255 2870 305 2885
rect 355 4055 405 4070
rect 355 2885 370 4055
rect 390 2885 405 4055
rect 355 2870 405 2885
rect 455 4055 505 4070
rect 455 2885 470 4055
rect 490 2885 505 4055
rect 455 2870 505 2885
rect 695 4055 745 4070
rect 695 2885 710 4055
rect 730 2885 745 4055
rect 695 2870 745 2885
rect 795 4055 845 4070
rect 795 2885 810 4055
rect 830 2885 845 4055
rect 795 2870 845 2885
rect 895 4055 945 4070
rect 895 2885 910 4055
rect 930 2885 945 4055
rect 895 2870 945 2885
rect 995 4055 1045 4070
rect 995 2885 1010 4055
rect 1030 2885 1045 4055
rect 995 2870 1045 2885
rect 1095 4055 1145 4070
rect 1095 2885 1110 4055
rect 1130 2885 1145 4055
rect 1095 2870 1145 2885
rect 1195 4055 1245 4070
rect 1195 2885 1210 4055
rect 1235 2885 1245 4055
rect 1195 2870 1245 2885
<< ndiffc >>
rect -35 1490 -10 2660
rect 70 1490 90 2660
rect 170 1490 190 2660
rect 270 1490 290 2660
rect 370 1490 390 2660
rect 470 1490 490 2660
rect 710 1490 730 2660
rect 810 1490 830 2660
rect 910 1490 930 2660
rect 1010 1490 1030 2660
rect 1110 1490 1130 2660
rect 1210 1490 1235 2660
rect -30 -30 -10 1140
rect 70 -30 90 1140
rect 170 -30 190 1140
rect 270 -30 290 1140
rect 370 -30 390 1140
rect 470 -30 490 1140
rect 710 -30 730 1140
rect 810 -30 830 1140
rect 910 -30 930 1140
rect 1010 -30 1030 1140
rect 1110 -30 1130 1140
rect 1210 -30 1230 1140
<< pdiffc >>
rect -35 2885 -10 4055
rect 70 2885 90 4055
rect 170 2885 190 4055
rect 270 2885 290 4055
rect 370 2885 390 4055
rect 470 2885 490 4055
rect 710 2885 730 4055
rect 810 2885 830 4055
rect 910 2885 930 4055
rect 1010 2885 1030 4055
rect 1110 2885 1130 4055
rect 1210 2885 1235 4055
<< psubdiff >>
rect -95 2660 -45 2675
rect -95 1490 -80 2660
rect -55 1490 -45 2660
rect -95 1475 -45 1490
rect 1245 2660 1295 2675
rect 1245 1490 1255 2660
rect 1280 1490 1295 2660
rect 1245 1475 1295 1490
rect -95 1140 -45 1155
rect -95 -30 -80 1140
rect -55 -30 -45 1140
rect -95 -45 -45 -30
rect 1245 1140 1295 1155
rect 1245 -30 1255 1140
rect 1280 -30 1295 1140
rect 1245 -45 1295 -30
<< nsubdiff >>
rect -95 4055 -45 4070
rect -95 2885 -80 4055
rect -55 2885 -45 4055
rect -95 2870 -45 2885
rect 1245 4055 1295 4070
rect 1245 2885 1255 4055
rect 1280 2885 1295 4055
rect 1245 2870 1295 2885
<< psubdiffcont >>
rect -80 1490 -55 2660
rect 1255 1490 1280 2660
rect -80 -30 -55 1140
rect 1255 -30 1280 1140
<< nsubdiffcont >>
rect -80 2885 -55 4055
rect 1255 2885 1280 4055
<< poly >>
rect 120 4215 160 4225
rect 120 4195 130 4215
rect 150 4195 160 4215
rect 120 4185 160 4195
rect 420 4215 460 4225
rect 420 4195 430 4215
rect 450 4195 460 4215
rect 420 4185 460 4195
rect 740 4215 780 4225
rect 740 4195 750 4215
rect 770 4195 780 4215
rect 740 4185 780 4195
rect 1040 4215 1080 4225
rect 1040 4195 1050 4215
rect 1070 4195 1080 4215
rect 1040 4185 1080 4195
rect 120 4130 135 4185
rect 430 4130 445 4185
rect 755 4130 770 4185
rect 1065 4130 1080 4185
rect 5 4115 55 4130
rect 5 4095 20 4115
rect 40 4095 55 4115
rect 5 4070 55 4095
rect 105 4115 155 4130
rect 105 4095 120 4115
rect 140 4095 155 4115
rect 105 4070 155 4095
rect 205 4115 255 4130
rect 205 4095 220 4115
rect 240 4095 255 4115
rect 205 4070 255 4095
rect 305 4115 355 4130
rect 305 4095 320 4115
rect 340 4095 355 4115
rect 305 4070 355 4095
rect 405 4115 455 4130
rect 405 4095 420 4115
rect 440 4095 455 4115
rect 405 4070 455 4095
rect 745 4115 795 4130
rect 745 4095 760 4115
rect 780 4095 795 4115
rect 745 4070 795 4095
rect 845 4115 895 4130
rect 845 4095 860 4115
rect 880 4095 895 4115
rect 845 4070 895 4095
rect 945 4115 995 4130
rect 945 4095 960 4115
rect 980 4095 995 4115
rect 945 4070 995 4095
rect 1045 4115 1095 4130
rect 1045 4095 1060 4115
rect 1080 4095 1095 4115
rect 1045 4070 1095 4095
rect 1145 4115 1195 4130
rect 1145 4095 1160 4115
rect 1180 4095 1195 4115
rect 1145 4070 1195 4095
rect 5 2845 55 2870
rect 105 2845 155 2870
rect 205 2845 255 2870
rect 305 2845 355 2870
rect 405 2845 455 2870
rect 745 2845 795 2870
rect 845 2845 895 2870
rect 945 2845 995 2870
rect 1045 2845 1095 2870
rect 1145 2845 1195 2870
rect 70 2815 1130 2820
rect 70 2795 80 2815
rect 105 2805 1095 2815
rect 105 2795 115 2805
rect 70 2790 115 2795
rect 5 2675 55 2700
rect 105 2675 155 2700
rect 205 2675 255 2700
rect 5 1455 55 1475
rect 5 1430 20 1455
rect 40 1430 55 1455
rect 5 1420 55 1430
rect 105 1455 155 1475
rect 105 1430 120 1455
rect 140 1430 155 1455
rect 105 1420 155 1430
rect 205 1420 255 1475
rect 215 1355 235 1420
rect 200 1350 245 1355
rect 200 1330 210 1350
rect 235 1330 245 1350
rect 200 1325 245 1330
rect 60 1220 105 1225
rect 60 1200 70 1220
rect 95 1210 105 1220
rect 325 1210 340 2805
rect 520 2770 565 2775
rect 520 2750 530 2770
rect 555 2750 565 2770
rect 520 2745 565 2750
rect 635 2770 680 2775
rect 635 2750 645 2770
rect 670 2750 680 2770
rect 635 2745 680 2750
rect 405 2675 455 2700
rect 405 1455 455 1475
rect 405 1430 420 1455
rect 440 1430 455 1455
rect 405 1420 455 1430
rect 415 1300 435 1420
rect 405 1295 450 1300
rect 405 1275 415 1295
rect 440 1275 450 1295
rect 405 1270 450 1275
rect 95 1200 340 1210
rect 60 1195 340 1200
rect 5 1155 55 1170
rect 105 1155 155 1170
rect 205 1155 255 1170
rect 305 1155 355 1170
rect 405 1155 455 1170
rect 520 1160 540 2745
rect 660 1160 680 2745
rect 745 2675 795 2700
rect 745 1455 795 1475
rect 745 1430 760 1455
rect 780 1430 795 1455
rect 745 1420 795 1430
rect 765 1300 785 1420
rect 750 1295 795 1300
rect 750 1275 760 1295
rect 785 1275 795 1295
rect 750 1270 795 1275
rect 860 1210 875 2805
rect 1085 2795 1095 2805
rect 1120 2795 1130 2815
rect 1085 2790 1130 2795
rect 945 2675 995 2700
rect 1045 2675 1095 2700
rect 1145 2675 1195 2700
rect 945 1420 995 1475
rect 1045 1455 1095 1475
rect 1045 1430 1060 1455
rect 1080 1430 1095 1455
rect 1045 1420 1095 1430
rect 1145 1455 1195 1475
rect 1145 1430 1160 1455
rect 1180 1430 1195 1455
rect 1145 1420 1195 1430
rect 965 1355 985 1420
rect 955 1350 1000 1355
rect 955 1330 965 1350
rect 990 1330 1000 1350
rect 955 1325 1000 1330
rect 1095 1220 1140 1225
rect 1095 1210 1105 1220
rect 860 1200 1105 1210
rect 1130 1200 1140 1220
rect 860 1195 1140 1200
rect 520 1155 565 1160
rect 520 1135 530 1155
rect 555 1135 565 1155
rect 520 1130 565 1135
rect 635 1155 680 1160
rect 745 1155 795 1170
rect 845 1155 895 1170
rect 945 1155 995 1170
rect 1045 1155 1095 1170
rect 1145 1155 1195 1170
rect 635 1135 645 1155
rect 670 1135 680 1155
rect 635 1130 680 1135
rect 5 -65 55 -45
rect 5 -90 20 -65
rect 40 -90 55 -65
rect 5 -100 55 -90
rect 105 -65 155 -45
rect 105 -90 120 -65
rect 140 -90 155 -65
rect 105 -100 155 -90
rect 205 -65 255 -45
rect 205 -90 220 -65
rect 240 -90 255 -65
rect 205 -100 255 -90
rect 305 -65 355 -45
rect 305 -90 320 -65
rect 340 -90 355 -65
rect 305 -100 355 -90
rect 405 -65 455 -45
rect 405 -90 420 -65
rect 440 -90 455 -65
rect 405 -100 455 -90
rect 480 -65 525 -60
rect 480 -85 490 -65
rect 515 -85 525 -65
rect 480 -90 525 -85
rect 675 -65 720 -60
rect 675 -85 685 -65
rect 710 -85 720 -65
rect 675 -90 720 -85
rect 320 -125 340 -100
rect 480 -125 500 -90
rect 320 -145 500 -125
rect 700 -125 720 -90
rect 745 -65 795 -45
rect 745 -90 760 -65
rect 780 -90 795 -65
rect 745 -100 795 -90
rect 845 -65 895 -45
rect 845 -90 860 -65
rect 880 -90 895 -65
rect 845 -100 895 -90
rect 945 -65 995 -45
rect 945 -90 960 -65
rect 980 -90 995 -65
rect 945 -100 995 -90
rect 1045 -65 1095 -45
rect 1045 -90 1060 -65
rect 1080 -90 1095 -65
rect 1045 -100 1095 -90
rect 1145 -65 1195 -45
rect 1145 -90 1160 -65
rect 1180 -90 1195 -65
rect 1145 -100 1195 -90
rect 860 -125 880 -100
rect 700 -145 880 -125
<< polycont >>
rect 130 4195 150 4215
rect 430 4195 450 4215
rect 750 4195 770 4215
rect 1050 4195 1070 4215
rect 20 4095 40 4115
rect 120 4095 140 4115
rect 220 4095 240 4115
rect 320 4095 340 4115
rect 420 4095 440 4115
rect 760 4095 780 4115
rect 860 4095 880 4115
rect 960 4095 980 4115
rect 1060 4095 1080 4115
rect 1160 4095 1180 4115
rect 80 2795 105 2815
rect 20 1430 40 1455
rect 120 1430 140 1455
rect 210 1330 235 1350
rect 70 1200 95 1220
rect 530 2750 555 2770
rect 645 2750 670 2770
rect 420 1430 440 1455
rect 415 1275 440 1295
rect 760 1430 780 1455
rect 760 1275 785 1295
rect 1095 2795 1120 2815
rect 1060 1430 1080 1455
rect 1160 1430 1180 1455
rect 965 1330 990 1350
rect 1105 1200 1130 1220
rect 530 1135 555 1155
rect 645 1135 670 1155
rect 20 -90 40 -65
rect 120 -90 140 -65
rect 220 -90 240 -65
rect 320 -90 340 -65
rect 420 -90 440 -65
rect 490 -85 515 -65
rect 685 -85 710 -65
rect 760 -90 780 -65
rect 860 -90 880 -65
rect 960 -90 980 -65
rect 1060 -90 1080 -65
rect 1160 -90 1180 -65
<< locali >>
rect 120 4215 160 4225
rect 120 4205 130 4215
rect -115 4195 130 4205
rect 150 4205 160 4215
rect 420 4215 460 4225
rect 420 4205 430 4215
rect 150 4195 430 4205
rect 450 4205 460 4215
rect 740 4215 780 4225
rect 740 4205 750 4215
rect 450 4195 750 4205
rect 770 4205 780 4215
rect 1040 4215 1080 4225
rect 1040 4205 1050 4215
rect 770 4195 1050 4205
rect 1070 4195 1080 4215
rect -115 4185 1080 4195
rect -115 4145 1080 4165
rect 230 4125 250 4145
rect 330 4125 350 4145
rect 850 4125 870 4145
rect 950 4125 970 4145
rect 10 4115 50 4125
rect 10 4105 20 4115
rect -20 4095 20 4105
rect 40 4095 50 4115
rect -20 4085 50 4095
rect 110 4115 150 4125
rect 110 4095 120 4115
rect 140 4095 150 4115
rect 110 4085 150 4095
rect 210 4115 250 4125
rect 210 4095 220 4115
rect 240 4095 250 4115
rect 210 4085 250 4095
rect 310 4115 350 4125
rect 310 4095 320 4115
rect 340 4095 350 4115
rect 310 4085 350 4095
rect 410 4115 450 4125
rect 410 4095 420 4115
rect 440 4095 450 4115
rect 410 4085 450 4095
rect 750 4115 790 4125
rect 750 4095 760 4115
rect 780 4095 790 4115
rect 750 4085 790 4095
rect 850 4115 890 4125
rect 850 4095 860 4115
rect 880 4095 890 4115
rect 850 4085 890 4095
rect 950 4115 990 4125
rect 950 4095 960 4115
rect 980 4095 990 4115
rect 950 4085 990 4095
rect 1050 4115 1090 4125
rect 1050 4095 1060 4115
rect 1080 4095 1090 4115
rect 1050 4085 1090 4095
rect 1150 4115 1190 4125
rect 1150 4095 1160 4115
rect 1180 4105 1190 4115
rect 1180 4095 1220 4105
rect 1150 4085 1220 4095
rect -20 4065 0 4085
rect 1200 4065 1220 4085
rect -90 4055 0 4065
rect -90 2885 -80 4055
rect -55 2885 -35 4055
rect -10 2885 0 4055
rect -90 2875 0 2885
rect 60 4055 100 4065
rect 60 2885 70 4055
rect 90 2885 100 4055
rect 60 2875 100 2885
rect 160 4055 200 4065
rect 160 2885 170 4055
rect 190 2885 200 4055
rect 160 2875 200 2885
rect 260 4055 300 4065
rect 260 2885 270 4055
rect 290 2885 300 4055
rect 260 2875 300 2885
rect 360 4055 400 4065
rect 360 2885 370 4055
rect 390 2885 400 4055
rect 360 2875 400 2885
rect 460 4055 500 4065
rect 460 2885 470 4055
rect 490 2895 500 4055
rect 700 4055 740 4065
rect 700 2895 710 4055
rect 490 2885 540 2895
rect 460 2875 540 2885
rect 70 2820 90 2875
rect 70 2815 115 2820
rect 70 2795 80 2815
rect 105 2795 115 2815
rect 70 2790 115 2795
rect 180 2750 200 2875
rect 360 2760 380 2875
rect 80 2730 200 2750
rect 280 2740 380 2760
rect 520 2775 540 2875
rect 660 2885 710 2895
rect 730 2885 740 4055
rect 660 2875 740 2885
rect 800 4055 840 4065
rect 800 2885 810 4055
rect 830 2885 840 4055
rect 800 2875 840 2885
rect 900 4055 940 4065
rect 900 2885 910 4055
rect 930 2885 940 4055
rect 900 2875 940 2885
rect 1000 4055 1040 4065
rect 1000 2885 1010 4055
rect 1030 2885 1040 4055
rect 1000 2875 1040 2885
rect 1100 4055 1140 4065
rect 1100 2885 1110 4055
rect 1130 2885 1140 4055
rect 1100 2875 1140 2885
rect 1200 4055 1290 4065
rect 1200 2885 1210 4055
rect 1235 2885 1255 4055
rect 1280 2885 1290 4055
rect 1200 2875 1290 2885
rect 660 2775 680 2875
rect 520 2770 565 2775
rect 520 2750 530 2770
rect 555 2750 565 2770
rect 520 2745 565 2750
rect 635 2770 680 2775
rect 635 2750 645 2770
rect 670 2750 680 2770
rect 635 2745 680 2750
rect 820 2760 840 2875
rect 820 2740 920 2760
rect 80 2670 100 2730
rect 280 2670 300 2740
rect 900 2670 920 2740
rect 1000 2750 1020 2875
rect 1110 2820 1130 2875
rect 1085 2815 1315 2820
rect 1085 2795 1095 2815
rect 1120 2800 1315 2815
rect 1120 2795 1130 2800
rect 1085 2790 1130 2795
rect 1000 2730 1120 2750
rect 1100 2670 1120 2730
rect -90 2660 0 2670
rect -90 1490 -80 2660
rect -55 1490 -35 2660
rect -10 1490 0 2660
rect -90 1480 0 1490
rect 60 2660 100 2670
rect 60 1490 70 2660
rect 90 1490 100 2660
rect 60 1480 100 1490
rect 160 2660 200 2670
rect 160 1490 170 2660
rect 190 1490 200 2660
rect 160 1480 200 1490
rect 260 2660 300 2670
rect 260 1490 270 2660
rect 290 1490 300 2660
rect 260 1480 300 1490
rect 360 2660 400 2670
rect 360 1490 370 2660
rect 390 1490 400 2660
rect 360 1480 400 1490
rect 460 2660 500 2670
rect 460 1490 470 2660
rect 490 1490 500 2660
rect 460 1480 500 1490
rect 700 2660 740 2670
rect 700 1490 710 2660
rect 730 1490 740 2660
rect 700 1480 740 1490
rect 800 2660 840 2670
rect 800 1490 810 2660
rect 830 1490 840 2660
rect 800 1480 840 1490
rect 900 2660 940 2670
rect 900 1490 910 2660
rect 930 1490 940 2660
rect 900 1480 940 1490
rect 1000 2660 1040 2670
rect 1000 1490 1010 2660
rect 1030 1490 1040 2660
rect 1000 1480 1040 1490
rect 1100 2660 1140 2670
rect 1100 1490 1110 2660
rect 1130 1490 1140 2660
rect 1100 1480 1140 1490
rect 1200 2660 1290 2670
rect 1200 1490 1210 2660
rect 1235 1490 1255 2660
rect 1280 1490 1290 2660
rect 1200 1480 1290 1490
rect -20 1460 0 1480
rect 180 1460 200 1480
rect 360 1460 380 1480
rect 820 1460 840 1480
rect 1000 1460 1020 1480
rect 1200 1460 1220 1480
rect -20 1455 50 1460
rect -20 1435 20 1455
rect 10 1430 20 1435
rect 40 1430 50 1455
rect 10 1425 50 1430
rect 110 1455 150 1460
rect 110 1430 120 1455
rect 140 1430 150 1455
rect 180 1440 380 1460
rect 410 1455 450 1460
rect 110 1425 150 1430
rect 410 1430 420 1455
rect 440 1430 450 1455
rect 410 1425 450 1430
rect 750 1455 790 1460
rect 750 1430 760 1455
rect 780 1430 790 1455
rect 820 1440 1020 1460
rect 1050 1455 1090 1460
rect 750 1425 790 1430
rect 1050 1430 1060 1455
rect 1080 1430 1090 1455
rect 1050 1425 1090 1430
rect 1150 1455 1220 1460
rect 1150 1430 1160 1455
rect 1180 1435 1220 1455
rect 1180 1430 1190 1435
rect 1150 1425 1190 1430
rect 120 1405 140 1425
rect 1060 1405 1080 1425
rect -115 1385 1080 1405
rect 200 1350 245 1355
rect 200 1340 210 1350
rect -115 1330 210 1340
rect 235 1340 245 1350
rect 955 1350 1000 1355
rect 955 1340 965 1350
rect 235 1330 965 1340
rect 990 1330 1000 1350
rect -115 1320 1000 1330
rect -115 1295 795 1300
rect -115 1280 415 1295
rect 405 1275 415 1280
rect 440 1280 760 1295
rect 440 1275 450 1280
rect 405 1270 450 1275
rect 750 1275 760 1280
rect 785 1275 795 1295
rect 750 1270 795 1275
rect 60 1220 105 1225
rect 60 1200 70 1220
rect 95 1200 105 1220
rect 60 1195 105 1200
rect 1095 1220 1140 1225
rect 1095 1200 1105 1220
rect 1130 1200 1140 1220
rect 1095 1195 1140 1200
rect 70 1150 90 1195
rect 520 1155 565 1160
rect 520 1150 530 1155
rect -90 1140 0 1150
rect -90 -30 -80 1140
rect -55 -30 -30 1140
rect -10 -30 0 1140
rect -90 -40 0 -30
rect 60 1140 100 1150
rect 60 -30 70 1140
rect 90 -30 100 1140
rect 60 -40 100 -30
rect 160 1140 200 1150
rect 160 -30 170 1140
rect 190 -30 200 1140
rect 160 -40 200 -30
rect 260 1140 300 1150
rect 260 -30 270 1140
rect 290 -30 300 1140
rect 260 -40 300 -30
rect 360 1140 400 1150
rect 360 -30 370 1140
rect 390 -30 400 1140
rect 360 -40 400 -30
rect 460 1140 530 1150
rect 460 -30 470 1140
rect 490 1135 530 1140
rect 555 1135 565 1155
rect 490 1130 565 1135
rect 635 1155 680 1160
rect 635 1135 645 1155
rect 670 1150 680 1155
rect 1110 1150 1130 1195
rect 670 1140 740 1150
rect 670 1135 710 1140
rect 635 1130 710 1135
rect 490 -30 500 1130
rect 460 -40 500 -30
rect -30 -65 -10 -40
rect 480 -60 500 -40
rect 700 -30 710 1130
rect 730 -30 740 1140
rect 700 -40 740 -30
rect 800 1140 840 1150
rect 800 -30 810 1140
rect 830 -30 840 1140
rect 800 -40 840 -30
rect 900 1140 940 1150
rect 900 -30 910 1140
rect 930 -30 940 1140
rect 900 -40 940 -30
rect 1000 1140 1040 1150
rect 1000 -30 1010 1140
rect 1030 -30 1040 1140
rect 1000 -40 1040 -30
rect 1100 1140 1140 1150
rect 1100 -30 1110 1140
rect 1130 -30 1140 1140
rect 1100 -40 1140 -30
rect 1200 1140 1290 1150
rect 1200 -30 1210 1140
rect 1230 -30 1255 1140
rect 1280 -30 1290 1140
rect 1200 -40 1290 -30
rect 700 -60 720 -40
rect 10 -65 50 -60
rect -30 -85 20 -65
rect 10 -90 20 -85
rect 40 -90 50 -65
rect 10 -95 50 -90
rect 110 -65 150 -60
rect 110 -90 120 -65
rect 140 -90 150 -65
rect 110 -95 150 -90
rect 210 -65 250 -60
rect 210 -90 220 -65
rect 240 -70 250 -65
rect 310 -65 350 -60
rect 310 -70 320 -65
rect 240 -90 320 -70
rect 340 -90 350 -65
rect 210 -95 250 -90
rect 310 -95 350 -90
rect 410 -65 450 -60
rect 410 -90 420 -65
rect 440 -90 450 -65
rect 480 -65 525 -60
rect 480 -85 490 -65
rect 515 -85 525 -65
rect 480 -90 525 -85
rect 675 -65 720 -60
rect 675 -85 685 -65
rect 710 -85 720 -65
rect 675 -90 720 -85
rect 750 -65 790 -60
rect 750 -90 760 -65
rect 780 -90 790 -65
rect 410 -95 450 -90
rect 750 -95 790 -90
rect 850 -65 890 -60
rect 850 -90 860 -65
rect 880 -70 890 -65
rect 950 -65 990 -60
rect 950 -70 960 -65
rect 880 -90 960 -70
rect 980 -90 990 -65
rect 850 -95 890 -90
rect 950 -95 990 -90
rect 1050 -65 1090 -60
rect 1050 -90 1060 -65
rect 1080 -90 1090 -65
rect 1050 -95 1090 -90
rect 1150 -65 1190 -60
rect 1210 -65 1230 -40
rect 1150 -90 1160 -65
rect 1180 -85 1230 -65
rect 1180 -90 1190 -85
rect 1150 -95 1190 -90
rect 120 -115 140 -95
rect 420 -115 440 -95
rect 760 -115 780 -95
rect 1060 -115 1080 -95
rect -115 -135 1080 -115
<< viali >>
rect -80 2885 -55 4055
rect -35 2885 -10 4055
rect 270 2885 290 4055
rect 910 2885 930 4055
rect 1210 2885 1235 4055
rect 1255 2885 1280 4055
rect -80 1490 -55 2660
rect -35 1490 -10 2660
rect 470 1490 490 2660
rect 710 1490 730 2660
rect 1210 1490 1235 2660
rect 1255 1490 1280 2660
rect -80 -30 -55 1140
rect -30 -30 -10 1140
rect 270 -30 290 1140
rect 910 -30 930 1140
rect 1210 -30 1230 1140
rect 1255 -30 1280 1140
<< metal1 >>
rect -115 4055 1315 4070
rect -115 2885 -80 4055
rect -55 2885 -35 4055
rect -10 2885 270 4055
rect 290 2885 910 4055
rect 930 2885 1210 4055
rect 1235 2885 1255 4055
rect 1280 2885 1315 4055
rect -115 2870 1315 2885
rect -115 2660 1315 2675
rect -115 1490 -80 2660
rect -55 1490 -35 2660
rect -10 1490 470 2660
rect 490 1490 710 2660
rect 730 1490 1210 2660
rect 1235 1490 1255 2660
rect 1280 1490 1315 2660
rect -115 1140 1315 1490
rect -115 -30 -80 1140
rect -55 -30 -30 1140
rect -10 -30 270 1140
rect 290 -30 910 1140
rect 930 -30 1210 1140
rect 1230 -30 1255 1140
rect 1280 -30 1315 1140
rect -115 -45 1315 -30
<< labels >>
rlabel locali -115 -125 -115 -125 7 VCN
port 1 w
rlabel locali -115 1290 -115 1290 7 VBN
port 2 w
rlabel locali -115 1330 -115 1330 7 V1
port 3 w
rlabel locali -115 1395 -115 1395 7 V2
port 4 w
rlabel locali -115 4155 -115 4155 7 VBP
port 5 w
rlabel locali -115 4195 -115 4195 7 VCP
port 6 w
rlabel locali 1315 2810 1315 2810 3 Vout
port 7 e
rlabel metal1 -115 1260 -115 1260 7 VN
port 8 w
rlabel metal1 -115 2885 -115 2885 7 VP
port 9 w
<< end >>
