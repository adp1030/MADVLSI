magic
tech sky130A
timestamp 1695859786
<< nwell >>
rect -240 545 585 1630
<< nmos >>
rect 215 365 230 465
rect 215 165 230 265
rect 10 -25 25 75
rect 75 -25 90 75
rect 365 -25 380 75
rect 430 -25 445 75
rect 215 -515 230 -115
<< pmos >>
rect 215 1170 230 1570
rect 10 980 25 1080
rect 75 980 90 1080
rect -130 780 -115 880
rect -130 580 -115 680
rect 365 975 380 1075
rect 430 975 445 1075
<< ndiff >>
rect 165 455 215 465
rect 165 375 180 455
rect 200 375 215 455
rect 165 365 215 375
rect 230 455 280 465
rect 230 375 245 455
rect 265 375 280 455
rect 230 365 280 375
rect 165 255 215 265
rect 165 175 180 255
rect 200 175 215 255
rect 165 165 215 175
rect 230 255 280 265
rect 230 175 245 255
rect 265 175 280 255
rect 230 165 280 175
rect -40 65 10 75
rect -40 -15 -25 65
rect -5 -15 10 65
rect -40 -25 10 -15
rect 25 65 75 75
rect 25 -15 40 65
rect 60 -15 75 65
rect 25 -25 75 -15
rect 90 65 140 75
rect 90 -15 105 65
rect 125 -15 140 65
rect 90 -25 140 -15
rect 315 65 365 75
rect 315 -15 330 65
rect 350 -15 365 65
rect 315 -25 365 -15
rect 380 65 430 75
rect 380 -15 395 65
rect 415 -15 430 65
rect 380 -25 430 -15
rect 445 65 495 75
rect 445 -15 460 65
rect 480 -15 495 65
rect 445 -25 495 -15
rect 165 -125 215 -115
rect 165 -205 180 -125
rect 200 -205 215 -125
rect 165 -515 215 -205
rect 230 -125 280 -115
rect 230 -205 245 -125
rect 265 -205 280 -125
rect 230 -515 280 -205
<< pdiff >>
rect 165 1260 215 1570
rect 165 1180 180 1260
rect 200 1180 215 1260
rect 165 1170 215 1180
rect 230 1260 280 1570
rect 230 1180 245 1260
rect 265 1180 280 1260
rect 230 1170 280 1180
rect -40 1070 10 1080
rect -40 990 -25 1070
rect -5 990 10 1070
rect -40 980 10 990
rect 25 1070 75 1080
rect 25 990 40 1070
rect 60 990 75 1070
rect 25 980 75 990
rect 90 1070 140 1080
rect 90 990 105 1070
rect 125 990 140 1070
rect 90 980 140 990
rect -180 870 -130 880
rect -180 790 -165 870
rect -145 790 -130 870
rect -180 780 -130 790
rect -115 870 -65 880
rect -115 790 -100 870
rect -80 790 -65 870
rect -115 780 -65 790
rect -180 670 -130 680
rect -180 590 -165 670
rect -145 590 -130 670
rect -180 580 -130 590
rect -115 670 -65 680
rect -115 590 -100 670
rect -80 590 -65 670
rect -115 580 -65 590
rect 315 1065 365 1075
rect 315 985 330 1065
rect 350 985 365 1065
rect 315 975 365 985
rect 380 1065 430 1075
rect 380 985 395 1065
rect 415 985 430 1065
rect 380 975 430 985
rect 445 1065 495 1075
rect 445 985 460 1065
rect 480 985 495 1065
rect 445 975 495 985
<< ndiffc >>
rect 180 375 200 455
rect 245 375 265 455
rect 180 175 200 255
rect 245 175 265 255
rect -25 -15 -5 65
rect 40 -15 60 65
rect 105 -15 125 65
rect 330 -15 350 65
rect 395 -15 415 65
rect 460 -15 480 65
rect 180 -205 200 -125
rect 245 -205 265 -125
<< pdiffc >>
rect 180 1180 200 1260
rect 245 1180 265 1260
rect -25 990 -5 1070
rect 40 990 60 1070
rect 105 990 125 1070
rect -165 790 -145 870
rect -100 790 -80 870
rect -165 590 -145 670
rect -100 590 -80 670
rect 330 985 350 1065
rect 395 985 415 1065
rect 460 985 480 1065
<< psubdiff >>
rect 415 -75 465 -65
rect 415 -155 430 -75
rect 450 -155 465 -75
rect 415 -165 465 -155
<< nsubdiff >>
rect 10 1205 60 1215
rect 10 1125 25 1205
rect 45 1125 60 1205
rect 10 1115 60 1125
<< psubdiffcont >>
rect 430 -155 450 -75
<< nsubdiffcont >>
rect 25 1125 45 1205
<< poly >>
rect 215 1570 230 1585
rect 10 1080 25 1095
rect 75 1080 90 1095
rect -110 960 -70 970
rect 10 960 25 980
rect -110 940 -100 960
rect -80 940 25 960
rect -110 930 -70 940
rect -130 880 -115 895
rect -130 680 -115 780
rect -130 -570 -115 580
rect 10 75 25 940
rect 75 315 90 980
rect 215 465 230 1170
rect 365 1075 380 1090
rect 430 1075 445 1090
rect 150 315 190 325
rect 75 295 160 315
rect 180 295 190 315
rect 75 75 90 295
rect 150 285 190 295
rect 215 265 230 365
rect 255 325 295 335
rect 365 325 380 975
rect 255 305 265 325
rect 285 305 380 325
rect 255 295 295 305
rect 10 -40 25 -25
rect 75 -40 90 -25
rect 215 -115 230 165
rect 365 75 380 305
rect 430 735 445 975
rect 510 735 550 745
rect 430 715 520 735
rect 540 715 550 735
rect 430 75 445 715
rect 510 705 550 715
rect 365 -40 380 -25
rect 430 -40 445 -25
rect 215 -570 230 -515
rect -130 -585 230 -570
rect 215 -610 230 -585
rect 205 -620 245 -610
rect 205 -640 215 -620
rect 235 -640 245 -620
rect 205 -650 245 -640
<< polycont >>
rect -100 940 -80 960
rect 160 295 180 315
rect 265 305 285 325
rect 520 715 540 735
rect 215 -640 235 -620
<< locali >>
rect 125 1595 370 1615
rect -110 1235 100 1255
rect -110 970 -90 1235
rect 15 1205 55 1210
rect 15 1125 25 1205
rect 45 1125 55 1205
rect 15 1120 55 1125
rect 35 1075 55 1120
rect 80 1115 100 1235
rect 125 1155 145 1595
rect 350 1275 370 1595
rect 170 1260 210 1265
rect 170 1180 180 1260
rect 200 1180 210 1260
rect 170 1175 210 1180
rect 235 1260 275 1265
rect 235 1180 245 1260
rect 265 1195 275 1260
rect 350 1255 470 1275
rect 265 1180 405 1195
rect 235 1175 405 1180
rect 125 1135 255 1155
rect 80 1095 195 1115
rect -35 1070 5 1075
rect -35 990 -25 1070
rect -5 990 5 1070
rect -35 985 5 990
rect 30 1070 70 1075
rect 30 990 40 1070
rect 60 990 70 1070
rect 30 985 70 990
rect 95 1070 135 1075
rect 95 990 105 1070
rect 125 990 135 1070
rect 95 985 135 990
rect -110 960 -70 970
rect -110 940 -100 960
rect -80 940 -70 960
rect -110 930 -70 940
rect -110 875 -90 930
rect -240 870 -135 875
rect -240 845 -165 870
rect -175 790 -165 845
rect -145 790 -135 870
rect -175 785 -135 790
rect -110 870 -70 875
rect -110 790 -100 870
rect -80 790 -70 870
rect -110 785 -70 790
rect -25 675 -5 985
rect -240 670 -135 675
rect -240 645 -165 670
rect -175 590 -165 645
rect -145 590 -135 670
rect -175 585 -135 590
rect -110 670 -5 675
rect -110 590 -100 670
rect -80 655 -5 670
rect -80 590 -70 655
rect -110 585 -70 590
rect -90 -535 -70 585
rect -25 70 -5 655
rect 105 420 125 985
rect 175 460 195 1095
rect 235 460 255 1135
rect 385 1070 405 1175
rect 450 1070 470 1255
rect 315 1065 360 1070
rect 315 985 330 1065
rect 350 985 360 1065
rect 315 980 360 985
rect 385 1065 425 1070
rect 385 985 395 1065
rect 415 985 425 1065
rect 385 980 425 985
rect 450 1065 490 1070
rect 450 985 460 1065
rect 480 1000 490 1065
rect 480 985 525 1000
rect 450 980 525 985
rect 170 455 210 460
rect 170 420 180 455
rect 105 400 180 420
rect 105 70 125 400
rect 170 375 180 400
rect 200 375 210 455
rect 170 370 210 375
rect 235 455 275 460
rect 235 375 245 455
rect 265 375 275 455
rect 235 370 275 375
rect 255 335 275 370
rect 255 325 295 335
rect 150 315 190 325
rect 150 295 160 315
rect 180 295 190 315
rect 255 305 265 325
rect 285 305 295 325
rect 255 295 295 305
rect 150 285 190 295
rect 170 260 190 285
rect 170 255 210 260
rect 170 175 180 255
rect 200 175 210 255
rect 170 170 210 175
rect 235 255 275 260
rect 235 175 245 255
rect 265 175 275 255
rect 235 170 275 175
rect 170 125 190 170
rect 170 105 235 125
rect -35 65 5 70
rect -35 -15 -25 65
rect -5 -15 5 65
rect -35 -20 5 -15
rect 30 65 70 70
rect 30 -15 40 65
rect 60 -15 70 65
rect 30 -20 70 -15
rect 95 65 140 70
rect 95 -15 105 65
rect 125 -15 140 65
rect 95 -20 140 -15
rect 50 -120 70 -20
rect 215 -40 235 105
rect 255 70 275 170
rect 330 70 350 980
rect 460 70 480 980
rect 505 875 525 980
rect 505 845 585 875
rect 510 735 550 745
rect 510 715 520 735
rect 540 715 550 735
rect 510 705 550 715
rect 510 675 530 705
rect 510 645 585 675
rect 255 65 360 70
rect 255 50 330 65
rect 320 -15 330 50
rect 350 -15 360 65
rect 320 -20 360 -15
rect 385 65 425 70
rect 385 -15 395 65
rect 415 -15 425 65
rect 385 -20 425 -15
rect 450 65 490 70
rect 450 -15 460 65
rect 480 -15 490 65
rect 450 -20 490 -15
rect 215 -60 320 -40
rect 50 -125 210 -120
rect 50 -140 180 -125
rect 170 -205 180 -140
rect 200 -205 210 -125
rect 170 -210 210 -205
rect 235 -125 275 -120
rect 235 -205 245 -125
rect 265 -205 275 -125
rect 235 -210 275 -205
rect 295 -535 320 -60
rect 340 -190 360 -20
rect 400 -70 420 -20
rect 400 -75 460 -70
rect 400 -100 430 -75
rect 420 -155 430 -100
rect 450 -155 460 -75
rect 420 -160 460 -155
rect 510 -190 530 645
rect 340 -210 530 -190
rect -90 -560 320 -535
rect 205 -620 245 -610
rect 205 -640 215 -620
rect 235 -640 245 -620
rect 205 -650 245 -640
<< viali >>
rect 25 1125 45 1205
rect 180 1180 200 1260
rect 40 990 60 1070
rect 395 -15 415 65
rect 245 -205 265 -125
rect 430 -155 450 -75
rect 215 -640 235 -620
<< metal1 >>
rect -240 1260 585 1615
rect -240 1205 180 1260
rect -240 1125 25 1205
rect 45 1180 180 1205
rect 200 1180 585 1260
rect 45 1125 585 1180
rect -240 1070 585 1125
rect -240 990 40 1070
rect 60 990 585 1070
rect -240 575 585 990
rect -240 65 585 470
rect -240 -15 395 65
rect 415 -15 585 65
rect -240 -75 585 -15
rect -240 -125 430 -75
rect -240 -205 245 -125
rect 265 -155 430 -125
rect 450 -155 585 -75
rect 265 -205 585 -155
rect -240 -560 585 -205
rect -240 -620 585 -610
rect -240 -640 215 -620
rect 235 -640 585 -620
rect -240 -650 585 -640
<< labels >>
rlabel locali -240 660 -240 660 7 Db
port 1 w
rlabel locali -240 860 -240 860 7 D
port 2 w
rlabel locali 585 860 585 860 3 Q
port 3 e
rlabel metal1 -240 1030 -240 1030 7 VP
port 5 w
rlabel metal1 -240 25 -240 25 7 VN
port 6 w
rlabel metal1 225 -650 225 -650 5 CLK
port 7 s
rlabel locali 585 660 585 660 3 Qb
port 4 e
<< end >>
