magic
tech sky130A
timestamp 1694201234
<< nwell >>
rect -440 45 -30 185
<< nmos >>
rect -320 -90 -305 10
rect -120 -90 -105 10
<< pmos >>
rect -320 65 -305 165
rect -120 65 -105 165
<< ndiff >>
rect -370 -5 -320 10
rect -370 -75 -355 -5
rect -335 -75 -320 -5
rect -370 -90 -320 -75
rect -305 -90 -120 10
rect -105 -5 -55 10
rect -105 -75 -90 -5
rect -70 -75 -55 -5
rect -105 -90 -55 -75
<< pdiff >>
rect -370 150 -320 165
rect -370 80 -355 150
rect -335 80 -320 150
rect -370 65 -320 80
rect -305 150 -255 165
rect -305 80 -290 150
rect -270 80 -255 150
rect -305 65 -255 80
rect -170 150 -120 165
rect -170 80 -155 150
rect -135 80 -120 150
rect -170 65 -120 80
rect -105 150 -55 165
rect -105 80 -90 150
rect -70 80 -55 150
rect -105 65 -55 80
<< ndiffc >>
rect -355 -75 -335 -5
rect -90 -75 -70 -5
<< pdiffc >>
rect -355 80 -335 150
rect -290 80 -270 150
rect -155 80 -135 150
rect -90 80 -70 150
<< psubdiff >>
rect -420 -5 -370 10
rect -420 -75 -405 -5
rect -385 -75 -370 -5
rect -420 -90 -370 -75
<< nsubdiff >>
rect -420 150 -370 165
rect -420 80 -405 150
rect -385 80 -370 150
rect -420 65 -370 80
rect -220 150 -170 165
rect -220 80 -205 150
rect -185 80 -170 150
rect -220 65 -170 80
<< psubdiffcont >>
rect -405 -75 -385 -5
<< nsubdiffcont >>
rect -405 80 -385 150
rect -205 80 -185 150
<< poly >>
rect -320 165 -305 180
rect -120 165 -105 180
rect -320 10 -305 65
rect -120 10 -105 65
rect -320 -105 -305 -90
rect -120 -105 -105 -90
rect -345 -115 -305 -105
rect -122 -106 -105 -105
rect -345 -135 -335 -115
rect -315 -135 -305 -115
rect -345 -145 -305 -135
rect -145 -115 -105 -106
rect -145 -135 -135 -115
rect -115 -135 -105 -115
rect -145 -145 -105 -135
<< polycont >>
rect -335 -135 -315 -115
rect -135 -135 -115 -115
<< locali >>
rect -290 200 -70 220
rect -290 160 -270 200
rect -90 160 -70 200
rect -415 150 -325 160
rect -415 80 -405 150
rect -385 80 -355 150
rect -335 80 -325 150
rect -415 70 -325 80
rect -300 150 -260 160
rect -300 80 -290 150
rect -270 80 -260 150
rect -300 70 -260 80
rect -215 150 -125 160
rect -215 80 -205 150
rect -185 80 -155 150
rect -135 80 -125 150
rect -215 70 -125 80
rect -100 150 -60 160
rect -100 80 -90 150
rect -70 80 -60 150
rect -100 70 -60 80
rect -80 5 -60 70
rect -415 -5 -325 5
rect -415 -75 -405 -5
rect -385 -75 -355 -5
rect -335 -75 -325 -5
rect -415 -85 -325 -75
rect -100 -5 -60 5
rect -100 -75 -90 -5
rect -70 -75 -60 -5
rect -100 -85 -60 -75
rect -80 -105 -60 -85
rect -345 -115 -305 -105
rect -122 -106 -105 -105
rect -345 -135 -335 -115
rect -315 -135 -305 -115
rect -345 -145 -305 -135
rect -145 -115 -105 -106
rect -145 -135 -135 -115
rect -115 -135 -105 -115
rect -80 -125 -30 -105
rect -145 -145 -105 -135
<< viali >>
rect -405 80 -385 150
rect -355 80 -335 150
rect -205 80 -185 150
rect -155 80 -135 150
rect -405 -75 -385 -5
rect -355 -75 -335 -5
<< metal1 >>
rect -440 150 -30 160
rect -440 80 -405 150
rect -385 80 -355 150
rect -335 80 -205 150
rect -185 80 -155 150
rect -135 80 -30 150
rect -440 70 -30 80
rect -440 -5 -29 5
rect -440 -75 -405 -5
rect -385 -75 -355 -5
rect -335 -75 -29 -5
rect -440 -85 -29 -75
<< labels >>
rlabel metal1 -440 115 -440 115 7 VP
port 4 w
rlabel metal1 -440 -35 -440 -35 7 VN
port 5 w
rlabel locali -30 -115 -30 -115 3 Y
port 3 e
rlabel locali -325 -145 -325 -145 5 B
port 2 s
rlabel locali -125 -145 -125 -145 5 A
port 1 s
rlabel ndiff -213 -88 -213 -88 5 VMID
<< end >>
