magic
tech sky130A
timestamp 1697606724
<< nwell >>
rect -120 2980 2650 5755
<< nmos >>
rect 0 1500 50 2700
rect 100 1500 150 2700
rect 340 1500 390 2700
rect 440 1500 490 2700
rect 540 1500 590 2700
rect 640 1500 690 2700
rect 820 1500 870 2700
rect 1060 1500 1110 2700
rect 0 0 50 1200
rect 100 0 150 1200
rect 280 0 330 1200
rect 460 0 510 1200
rect 640 0 690 1200
rect 820 0 870 1200
rect 1060 0 1110 1200
rect 1420 1500 1470 2700
rect 1660 1500 1710 2700
rect 1840 1500 1890 2700
rect 1940 1500 1990 2700
rect 2040 1500 2090 2700
rect 2140 1500 2190 2700
rect 2380 1500 2430 2700
rect 2480 1500 2530 2700
rect 1420 0 1470 1200
rect 1660 0 1710 1200
rect 1840 0 1890 1200
rect 2020 0 2070 1200
rect 2200 0 2250 1200
rect 2380 0 2430 1200
rect 2480 0 2530 1200
<< pmos >>
rect 0 4500 50 5700
rect 100 4500 150 5700
rect 340 4500 390 5700
rect 440 4500 490 5700
rect 540 4500 590 5700
rect 640 4500 690 5700
rect 1060 4500 1110 5700
rect 1420 4500 1470 5700
rect 1840 4500 1890 5700
rect 1940 4500 1990 5700
rect 2040 4500 2090 5700
rect 2140 4500 2190 5700
rect 2380 4500 2430 5700
rect 2480 4500 2530 5700
rect 0 3000 50 4200
rect 100 3000 150 4200
rect 280 3000 330 4200
rect 460 3000 510 4200
rect 640 3000 690 4200
rect 820 3000 870 4200
rect 1060 3000 1110 4200
rect 1420 3000 1470 4200
rect 1660 3000 1710 4200
rect 1840 3000 1890 4200
rect 2020 3000 2070 4200
rect 2200 3000 2250 4200
rect 2380 3000 2430 4200
rect 2480 3000 2530 4200
<< ndiff >>
rect -50 2685 0 2700
rect -50 1515 -35 2685
rect -15 1515 0 2685
rect -50 1500 0 1515
rect 50 2685 100 2700
rect 50 1515 65 2685
rect 85 1515 100 2685
rect 50 1500 100 1515
rect 150 2685 200 2700
rect 150 1515 165 2685
rect 185 1515 200 2685
rect 150 1500 200 1515
rect 290 2685 340 2700
rect 290 1515 305 2685
rect 325 1515 340 2685
rect 290 1500 340 1515
rect 390 2685 440 2700
rect 390 1515 405 2685
rect 425 1515 440 2685
rect 390 1500 440 1515
rect 490 2685 540 2700
rect 490 1515 505 2685
rect 525 1515 540 2685
rect 490 1500 540 1515
rect 590 2685 640 2700
rect 590 1515 605 2685
rect 625 1515 640 2685
rect 590 1500 640 1515
rect 690 2685 740 2700
rect 690 1515 705 2685
rect 725 1515 740 2685
rect 690 1500 740 1515
rect 770 2685 820 2700
rect 770 1515 785 2685
rect 805 1515 820 2685
rect 770 1500 820 1515
rect 870 2685 920 2700
rect 870 1515 885 2685
rect 905 1515 920 2685
rect 870 1500 920 1515
rect 1010 2685 1060 2700
rect 1010 1515 1025 2685
rect 1045 1515 1060 2685
rect 1010 1500 1060 1515
rect 1110 2685 1160 2700
rect 1110 1515 1125 2685
rect 1145 1515 1160 2685
rect 1370 2685 1420 2700
rect 1110 1500 1160 1515
rect -50 1185 0 1200
rect -50 15 -35 1185
rect -15 15 0 1185
rect -50 0 0 15
rect 50 1185 100 1200
rect 50 15 65 1185
rect 85 15 100 1185
rect 50 0 100 15
rect 150 1185 200 1200
rect 150 15 165 1185
rect 185 15 200 1185
rect 150 0 200 15
rect 230 1185 280 1200
rect 230 15 245 1185
rect 265 15 280 1185
rect 230 0 280 15
rect 330 1185 380 1200
rect 330 15 345 1185
rect 365 15 380 1185
rect 330 0 380 15
rect 410 1185 460 1200
rect 410 15 425 1185
rect 445 15 460 1185
rect 410 0 460 15
rect 510 1185 560 1200
rect 510 15 525 1185
rect 545 15 560 1185
rect 510 0 560 15
rect 590 1185 640 1200
rect 590 15 605 1185
rect 625 15 640 1185
rect 590 0 640 15
rect 690 1185 740 1200
rect 690 15 705 1185
rect 725 15 740 1185
rect 690 0 740 15
rect 770 1185 820 1200
rect 770 15 785 1185
rect 805 15 820 1185
rect 770 0 820 15
rect 870 1185 920 1200
rect 870 15 885 1185
rect 905 15 920 1185
rect 870 0 920 15
rect 1010 1185 1060 1200
rect 1010 15 1025 1185
rect 1045 15 1060 1185
rect 1010 0 1060 15
rect 1110 1185 1160 1200
rect 1110 15 1125 1185
rect 1145 15 1160 1185
rect 1370 1515 1385 2685
rect 1405 1515 1420 2685
rect 1370 1500 1420 1515
rect 1470 2685 1520 2700
rect 1470 1515 1485 2685
rect 1505 1515 1520 2685
rect 1470 1500 1520 1515
rect 1610 2685 1660 2700
rect 1610 1515 1625 2685
rect 1645 1515 1660 2685
rect 1610 1500 1660 1515
rect 1710 2685 1760 2700
rect 1710 1515 1725 2685
rect 1745 1515 1760 2685
rect 1710 1500 1760 1515
rect 1790 2685 1840 2700
rect 1790 1515 1805 2685
rect 1825 1515 1840 2685
rect 1790 1500 1840 1515
rect 1890 2685 1940 2700
rect 1890 1515 1905 2685
rect 1925 1515 1940 2685
rect 1890 1500 1940 1515
rect 1990 2685 2040 2700
rect 1990 1515 2005 2685
rect 2025 1515 2040 2685
rect 1990 1500 2040 1515
rect 2090 2685 2140 2700
rect 2090 1515 2105 2685
rect 2125 1515 2140 2685
rect 2090 1500 2140 1515
rect 2190 2685 2240 2700
rect 2190 1515 2205 2685
rect 2225 1515 2240 2685
rect 2190 1500 2240 1515
rect 2330 2685 2380 2700
rect 2330 1515 2345 2685
rect 2365 1515 2380 2685
rect 2330 1500 2380 1515
rect 2430 2685 2480 2700
rect 2430 1515 2445 2685
rect 2465 1515 2480 2685
rect 2430 1500 2480 1515
rect 2530 2685 2580 2700
rect 2530 1515 2545 2685
rect 2565 1515 2580 2685
rect 2530 1500 2580 1515
rect 1370 1185 1420 1200
rect 1110 0 1160 15
rect 1370 15 1385 1185
rect 1405 15 1420 1185
rect 1370 0 1420 15
rect 1470 1185 1520 1200
rect 1470 15 1485 1185
rect 1505 15 1520 1185
rect 1470 0 1520 15
rect 1610 1185 1660 1200
rect 1610 15 1625 1185
rect 1645 15 1660 1185
rect 1610 0 1660 15
rect 1710 1185 1760 1200
rect 1710 15 1725 1185
rect 1745 15 1760 1185
rect 1710 0 1760 15
rect 1790 1185 1840 1200
rect 1790 15 1805 1185
rect 1825 15 1840 1185
rect 1790 0 1840 15
rect 1890 1185 1940 1200
rect 1890 15 1905 1185
rect 1925 15 1940 1185
rect 1890 0 1940 15
rect 1970 1185 2020 1200
rect 1970 15 1985 1185
rect 2005 15 2020 1185
rect 1970 0 2020 15
rect 2070 1185 2120 1200
rect 2070 15 2085 1185
rect 2105 15 2120 1185
rect 2070 0 2120 15
rect 2150 1185 2200 1200
rect 2150 15 2165 1185
rect 2185 15 2200 1185
rect 2150 0 2200 15
rect 2250 1185 2300 1200
rect 2250 15 2265 1185
rect 2285 15 2300 1185
rect 2250 0 2300 15
rect 2330 1185 2380 1200
rect 2330 15 2345 1185
rect 2365 15 2380 1185
rect 2330 0 2380 15
rect 2430 1185 2480 1200
rect 2430 15 2445 1185
rect 2465 15 2480 1185
rect 2430 0 2480 15
rect 2530 1185 2580 1200
rect 2530 15 2545 1185
rect 2565 15 2580 1185
rect 2530 0 2580 15
<< pdiff >>
rect -50 5685 0 5700
rect -50 4515 -35 5685
rect -15 4515 0 5685
rect -50 4500 0 4515
rect 50 5685 100 5700
rect 50 4515 65 5685
rect 85 4515 100 5685
rect 50 4500 100 4515
rect 150 5685 200 5700
rect 150 4515 165 5685
rect 185 4515 200 5685
rect 150 4500 200 4515
rect 290 5685 340 5700
rect 290 4515 305 5685
rect 325 4515 340 5685
rect 290 4500 340 4515
rect 390 5685 440 5700
rect 390 4515 405 5685
rect 425 4515 440 5685
rect 390 4500 440 4515
rect 490 5685 540 5700
rect 490 4515 505 5685
rect 525 4515 540 5685
rect 490 4500 540 4515
rect 590 5685 640 5700
rect 590 4515 605 5685
rect 625 4515 640 5685
rect 590 4500 640 4515
rect 690 5685 740 5700
rect 690 4515 705 5685
rect 725 4515 740 5685
rect 690 4500 740 4515
rect 1010 5685 1060 5700
rect 1010 4515 1025 5685
rect 1045 4515 1060 5685
rect 1010 4500 1060 4515
rect 1110 5685 1160 5700
rect 1110 4515 1125 5685
rect 1145 4515 1160 5685
rect 1110 4500 1160 4515
rect 1370 5685 1420 5700
rect 1370 4515 1385 5685
rect 1405 4515 1420 5685
rect 1370 4500 1420 4515
rect 1470 5685 1520 5700
rect 1470 4515 1485 5685
rect 1505 4515 1520 5685
rect 1470 4500 1520 4515
rect 1790 5685 1840 5700
rect 1790 4515 1805 5685
rect 1825 4515 1840 5685
rect 1790 4500 1840 4515
rect 1890 5685 1940 5700
rect 1890 4515 1905 5685
rect 1925 4515 1940 5685
rect 1890 4500 1940 4515
rect 1990 5685 2040 5700
rect 1990 4515 2005 5685
rect 2025 4515 2040 5685
rect 1990 4500 2040 4515
rect 2090 5685 2140 5700
rect 2090 4515 2105 5685
rect 2125 4515 2140 5685
rect 2090 4500 2140 4515
rect 2190 5685 2240 5700
rect 2190 4515 2205 5685
rect 2225 4515 2240 5685
rect 2190 4500 2240 4515
rect 2330 5685 2380 5700
rect 2330 4515 2345 5685
rect 2365 4515 2380 5685
rect 2330 4500 2380 4515
rect 2430 5685 2480 5700
rect 2430 4515 2445 5685
rect 2465 4515 2480 5685
rect 2430 4500 2480 4515
rect 2530 5685 2580 5700
rect 2530 4515 2545 5685
rect 2565 4515 2580 5685
rect 2530 4500 2580 4515
rect -50 4185 0 4200
rect -50 3015 -35 4185
rect -15 3015 0 4185
rect -50 3000 0 3015
rect 50 4185 100 4200
rect 50 3015 65 4185
rect 85 3015 100 4185
rect 50 3000 100 3015
rect 150 4185 200 4200
rect 150 3015 165 4185
rect 185 3015 200 4185
rect 150 3000 200 3015
rect 230 4185 280 4200
rect 230 3015 245 4185
rect 265 3015 280 4185
rect 230 3000 280 3015
rect 330 4185 380 4200
rect 330 3015 345 4185
rect 365 3015 380 4185
rect 330 3000 380 3015
rect 410 4185 460 4200
rect 410 3015 425 4185
rect 445 3015 460 4185
rect 410 3000 460 3015
rect 510 4185 560 4200
rect 510 3015 525 4185
rect 545 3015 560 4185
rect 510 3000 560 3015
rect 590 4185 640 4200
rect 590 3015 605 4185
rect 625 3015 640 4185
rect 590 3000 640 3015
rect 690 4185 740 4200
rect 690 3015 705 4185
rect 725 3015 740 4185
rect 690 3000 740 3015
rect 770 4185 820 4200
rect 770 3015 785 4185
rect 805 3015 820 4185
rect 770 3000 820 3015
rect 870 4185 920 4200
rect 870 3015 885 4185
rect 905 3015 920 4185
rect 870 3000 920 3015
rect 1010 4185 1060 4200
rect 1010 3015 1025 4185
rect 1045 3015 1060 4185
rect 1010 3000 1060 3015
rect 1110 4185 1160 4200
rect 1110 3015 1125 4185
rect 1145 3015 1160 4185
rect 1110 3000 1160 3015
rect 1370 4185 1420 4200
rect 1370 3015 1385 4185
rect 1405 3015 1420 4185
rect 1370 3000 1420 3015
rect 1470 4185 1520 4200
rect 1470 3015 1485 4185
rect 1505 3015 1520 4185
rect 1470 3000 1520 3015
rect 1610 4185 1660 4200
rect 1610 3015 1625 4185
rect 1645 3015 1660 4185
rect 1610 3000 1660 3015
rect 1710 4185 1760 4200
rect 1710 3015 1725 4185
rect 1745 3015 1760 4185
rect 1710 3000 1760 3015
rect 1790 4185 1840 4200
rect 1790 3015 1805 4185
rect 1825 3015 1840 4185
rect 1790 3000 1840 3015
rect 1890 4185 1940 4200
rect 1890 3015 1905 4185
rect 1925 3015 1940 4185
rect 1890 3000 1940 3015
rect 1970 4185 2020 4200
rect 1970 3015 1985 4185
rect 2005 3015 2020 4185
rect 1970 3000 2020 3015
rect 2070 4185 2120 4200
rect 2070 3015 2085 4185
rect 2105 3015 2120 4185
rect 2070 3000 2120 3015
rect 2150 4185 2200 4200
rect 2150 3015 2165 4185
rect 2185 3015 2200 4185
rect 2150 3000 2200 3015
rect 2250 4185 2300 4200
rect 2250 3015 2265 4185
rect 2285 3015 2300 4185
rect 2250 3000 2300 3015
rect 2330 4185 2380 4200
rect 2330 3015 2345 4185
rect 2365 3015 2380 4185
rect 2330 3000 2380 3015
rect 2430 4185 2480 4200
rect 2430 3015 2445 4185
rect 2465 3015 2480 4185
rect 2430 3000 2480 3015
rect 2530 4185 2580 4200
rect 2530 3015 2545 4185
rect 2565 3015 2580 4185
rect 2530 3000 2580 3015
<< ndiffc >>
rect -35 1515 -15 2685
rect 65 1515 85 2685
rect 165 1515 185 2685
rect 305 1515 325 2685
rect 405 1515 425 2685
rect 505 1515 525 2685
rect 605 1515 625 2685
rect 705 1515 725 2685
rect 785 1515 805 2685
rect 885 1515 905 2685
rect 1025 1515 1045 2685
rect 1125 1515 1145 2685
rect -35 15 -15 1185
rect 65 15 85 1185
rect 165 15 185 1185
rect 245 15 265 1185
rect 345 15 365 1185
rect 425 15 445 1185
rect 525 15 545 1185
rect 605 15 625 1185
rect 705 15 725 1185
rect 785 15 805 1185
rect 885 15 905 1185
rect 1025 15 1045 1185
rect 1125 15 1145 1185
rect 1385 1515 1405 2685
rect 1485 1515 1505 2685
rect 1625 1515 1645 2685
rect 1725 1515 1745 2685
rect 1805 1515 1825 2685
rect 1905 1515 1925 2685
rect 2005 1515 2025 2685
rect 2105 1515 2125 2685
rect 2205 1515 2225 2685
rect 2345 1515 2365 2685
rect 2445 1515 2465 2685
rect 2545 1515 2565 2685
rect 1385 15 1405 1185
rect 1485 15 1505 1185
rect 1625 15 1645 1185
rect 1725 15 1745 1185
rect 1805 15 1825 1185
rect 1905 15 1925 1185
rect 1985 15 2005 1185
rect 2085 15 2105 1185
rect 2165 15 2185 1185
rect 2265 15 2285 1185
rect 2345 15 2365 1185
rect 2445 15 2465 1185
rect 2545 15 2565 1185
<< pdiffc >>
rect -35 4515 -15 5685
rect 65 4515 85 5685
rect 165 4515 185 5685
rect 305 4515 325 5685
rect 405 4515 425 5685
rect 505 4515 525 5685
rect 605 4515 625 5685
rect 705 4515 725 5685
rect 1025 4515 1045 5685
rect 1125 4515 1145 5685
rect 1385 4515 1405 5685
rect 1485 4515 1505 5685
rect 1805 4515 1825 5685
rect 1905 4515 1925 5685
rect 2005 4515 2025 5685
rect 2105 4515 2125 5685
rect 2205 4515 2225 5685
rect 2345 4515 2365 5685
rect 2445 4515 2465 5685
rect 2545 4515 2565 5685
rect -35 3015 -15 4185
rect 65 3015 85 4185
rect 165 3015 185 4185
rect 245 3015 265 4185
rect 345 3015 365 4185
rect 425 3015 445 4185
rect 525 3015 545 4185
rect 605 3015 625 4185
rect 705 3015 725 4185
rect 785 3015 805 4185
rect 885 3015 905 4185
rect 1025 3015 1045 4185
rect 1125 3015 1145 4185
rect 1385 3015 1405 4185
rect 1485 3015 1505 4185
rect 1625 3015 1645 4185
rect 1725 3015 1745 4185
rect 1805 3015 1825 4185
rect 1905 3015 1925 4185
rect 1985 3015 2005 4185
rect 2085 3015 2105 4185
rect 2165 3015 2185 4185
rect 2265 3015 2285 4185
rect 2345 3015 2365 4185
rect 2445 3015 2465 4185
rect 2545 3015 2565 4185
<< psubdiff >>
rect -100 2685 -50 2700
rect -100 1515 -85 2685
rect -60 1515 -50 2685
rect -100 1500 -50 1515
rect -100 1185 -50 1200
rect -100 15 -85 1185
rect -60 15 -50 1185
rect -100 0 -50 15
rect 2580 2685 2630 2700
rect 2580 1515 2590 2685
rect 2615 1515 2630 2685
rect 2580 1500 2630 1515
rect 2580 1185 2630 1200
rect 2580 15 2590 1185
rect 2615 15 2630 1185
rect 2580 0 2630 15
<< nsubdiff >>
rect -100 5685 -50 5700
rect -100 4515 -85 5685
rect -60 4515 -50 5685
rect -100 4500 -50 4515
rect 2580 5685 2630 5700
rect 2580 4515 2590 5685
rect 2615 4515 2630 5685
rect 2580 4500 2630 4515
rect -100 4185 -50 4200
rect -100 3015 -85 4185
rect -60 3015 -50 4185
rect -100 3000 -50 3015
rect 2580 4185 2630 4200
rect 2580 3015 2590 4185
rect 2615 3015 2630 4185
rect 2580 3000 2630 3015
<< psubdiffcont >>
rect -85 1515 -60 2685
rect -85 15 -60 1185
rect 2590 1515 2615 2685
rect 2590 15 2615 1185
<< nsubdiffcont >>
rect -85 4515 -60 5685
rect 2590 4515 2615 5685
rect -85 3015 -60 4185
rect 2590 3015 2615 4185
<< poly >>
rect 1280 5765 1320 5770
rect 1280 5755 1290 5765
rect 0 5745 50 5755
rect 0 5725 15 5745
rect 35 5725 50 5745
rect 0 5700 50 5725
rect 100 5700 150 5755
rect 340 5745 1290 5755
rect 1310 5755 1320 5765
rect 1310 5745 2190 5755
rect 340 5725 965 5745
rect 985 5725 1075 5745
rect 1095 5740 1435 5745
rect 1095 5725 1180 5740
rect 340 5715 1180 5725
rect 1350 5725 1435 5740
rect 1455 5725 1545 5745
rect 1565 5725 2190 5745
rect 1350 5715 2190 5725
rect 340 5700 390 5715
rect 440 5700 490 5715
rect 540 5700 590 5715
rect 640 5700 690 5715
rect 1060 5700 1110 5715
rect 1420 5700 1470 5715
rect 1840 5700 1890 5715
rect 1940 5700 1990 5715
rect 2040 5700 2090 5715
rect 2140 5700 2190 5715
rect 2380 5700 2430 5755
rect 2480 5745 2530 5755
rect 2480 5725 2495 5745
rect 2515 5725 2530 5745
rect 2480 5700 2530 5725
rect 0 4485 50 4500
rect 100 4255 150 4500
rect 340 4485 390 4500
rect 440 4485 490 4500
rect 540 4485 590 4500
rect 640 4485 690 4500
rect 1060 4475 1110 4500
rect 1060 4455 1075 4475
rect 1095 4455 1110 4475
rect 1060 4445 1110 4455
rect 1420 4475 1470 4500
rect 1840 4485 1890 4500
rect 1940 4485 1990 4500
rect 2040 4485 2090 4500
rect 2140 4485 2190 4500
rect 1420 4455 1435 4475
rect 1455 4455 1470 4475
rect 1420 4445 1470 4455
rect 1200 4340 1240 4345
rect 1200 4330 1210 4340
rect 835 4320 1210 4330
rect 1230 4330 1240 4340
rect 1230 4320 1695 4330
rect 835 4315 1695 4320
rect 835 4255 855 4315
rect 1675 4255 1695 4315
rect 2380 4255 2430 4500
rect 2480 4485 2530 4500
rect 0 4245 50 4255
rect 0 4225 15 4245
rect 35 4225 50 4245
rect 0 4200 50 4225
rect 100 4245 690 4255
rect 100 4225 115 4245
rect 135 4225 295 4245
rect 315 4225 475 4245
rect 495 4225 655 4245
rect 675 4225 690 4245
rect 100 4215 690 4225
rect 100 4200 150 4215
rect 280 4200 330 4215
rect 460 4200 510 4215
rect 640 4200 690 4215
rect 820 4245 870 4255
rect 820 4225 835 4245
rect 855 4225 870 4245
rect 820 4200 870 4225
rect 1060 4245 1110 4255
rect 1060 4225 1075 4245
rect 1095 4225 1110 4245
rect 1060 4200 1110 4225
rect 1420 4245 1470 4255
rect 1420 4225 1435 4245
rect 1455 4225 1470 4245
rect 1420 4200 1470 4225
rect 1660 4245 1710 4255
rect 1660 4225 1675 4245
rect 1695 4225 1710 4245
rect 1660 4200 1710 4225
rect 1840 4245 2430 4255
rect 1840 4225 1855 4245
rect 1875 4225 2035 4245
rect 2055 4225 2215 4245
rect 2235 4225 2395 4245
rect 2415 4225 2430 4245
rect 1840 4215 2430 4225
rect 1840 4200 1890 4215
rect 2020 4200 2070 4215
rect 2200 4200 2250 4215
rect 2380 4200 2430 4215
rect 2480 4245 2530 4255
rect 2480 4225 2495 4245
rect 2515 4225 2530 4245
rect 2480 4200 2530 4225
rect 0 2985 50 3000
rect 100 2985 150 3000
rect 280 2985 330 3000
rect 460 2985 510 3000
rect 640 2985 690 3000
rect 820 2985 870 3000
rect 1060 2985 1110 3000
rect 1420 2985 1470 3000
rect 1660 2985 1710 3000
rect 1840 2985 1890 3000
rect 2020 2985 2070 3000
rect 2200 2985 2250 3000
rect 2380 2985 2430 3000
rect 2480 2985 2530 3000
rect 0 2745 50 2755
rect 0 2720 15 2745
rect 35 2720 50 2745
rect 0 2700 50 2720
rect 100 2745 1110 2755
rect 100 2720 115 2745
rect 135 2725 1110 2745
rect 1420 2745 2430 2755
rect 1420 2725 2395 2745
rect 135 2720 2395 2725
rect 2415 2720 2430 2745
rect 100 2715 2430 2720
rect 100 2700 150 2715
rect 340 2700 390 2715
rect 440 2700 490 2715
rect 540 2700 590 2715
rect 640 2700 690 2715
rect 820 2700 870 2715
rect 1060 2710 1470 2715
rect 1060 2700 1110 2710
rect 1420 2700 1470 2710
rect 1660 2700 1710 2715
rect 1840 2700 1890 2715
rect 1940 2700 1990 2715
rect 2040 2700 2090 2715
rect 2140 2700 2190 2715
rect 2380 2700 2430 2715
rect 2480 2745 2530 2755
rect 2480 2720 2495 2745
rect 2515 2720 2530 2745
rect 2480 2700 2530 2720
rect 1175 1950 1220 1955
rect 1175 1930 1185 1950
rect 1210 1930 1220 1950
rect 1175 1925 1220 1930
rect 1310 1950 1355 1955
rect 1310 1930 1320 1950
rect 1345 1930 1355 1950
rect 1310 1925 1355 1930
rect 0 1485 50 1500
rect 100 1485 150 1500
rect 340 1485 390 1500
rect 440 1485 490 1500
rect 540 1485 590 1500
rect 640 1485 690 1500
rect 820 1485 870 1500
rect 1060 1485 1110 1500
rect 1175 1255 1190 1925
rect 1270 1295 1310 1305
rect 1270 1275 1280 1295
rect 1300 1275 1310 1295
rect 1270 1265 1310 1275
rect 0 1245 50 1255
rect 0 1220 15 1245
rect 35 1220 50 1245
rect 0 1200 50 1220
rect 100 1245 870 1255
rect 100 1220 115 1245
rect 135 1220 295 1245
rect 315 1220 475 1245
rect 495 1220 655 1245
rect 675 1220 835 1245
rect 855 1220 870 1245
rect 100 1215 870 1220
rect 100 1200 150 1215
rect 280 1200 330 1215
rect 460 1200 510 1215
rect 640 1200 690 1215
rect 820 1200 870 1215
rect 1060 1245 1190 1255
rect 1060 1220 1075 1245
rect 1095 1240 1190 1245
rect 1095 1220 1110 1240
rect 1060 1200 1110 1220
rect 1280 1145 1295 1265
rect 1340 1255 1355 1925
rect 1420 1485 1470 1500
rect 1660 1485 1710 1500
rect 1840 1485 1890 1500
rect 1940 1485 1990 1500
rect 2040 1485 2090 1500
rect 2140 1485 2190 1500
rect 2380 1485 2430 1500
rect 2480 1485 2530 1500
rect 1340 1245 1470 1255
rect 1340 1240 1435 1245
rect 1420 1220 1435 1240
rect 1455 1220 1470 1245
rect 1420 1200 1470 1220
rect 1660 1245 2430 1255
rect 1660 1220 1675 1245
rect 1695 1220 1855 1245
rect 1875 1220 2035 1245
rect 2055 1220 2215 1245
rect 2235 1220 2395 1245
rect 2415 1220 2430 1245
rect 1660 1215 2430 1220
rect 1660 1200 1710 1215
rect 1840 1200 1890 1215
rect 2020 1200 2070 1215
rect 2200 1200 2250 1215
rect 2380 1200 2430 1215
rect 2480 1245 2530 1255
rect 2480 1220 2495 1245
rect 2515 1220 2530 1245
rect 2480 1200 2530 1220
rect 1270 1135 1310 1145
rect 1270 1115 1280 1135
rect 1300 1115 1310 1135
rect 1270 1105 1310 1115
rect 0 -15 50 0
rect 100 -15 150 0
rect 280 -15 330 0
rect 460 -15 510 0
rect 640 -15 690 0
rect 820 -15 870 0
rect 1060 -15 1110 0
rect 1420 -15 1470 0
rect 1660 -15 1710 0
rect 1840 -15 1890 0
rect 2020 -15 2070 0
rect 2200 -15 2250 0
rect 2380 -15 2430 0
rect 2480 -15 2530 0
<< polycont >>
rect 15 5725 35 5745
rect 1290 5745 1310 5765
rect 965 5725 985 5745
rect 1075 5725 1095 5745
rect 1435 5725 1455 5745
rect 1545 5725 1565 5745
rect 2495 5725 2515 5745
rect 1075 4455 1095 4475
rect 1435 4455 1455 4475
rect 1210 4320 1230 4340
rect 15 4225 35 4245
rect 115 4225 135 4245
rect 295 4225 315 4245
rect 475 4225 495 4245
rect 655 4225 675 4245
rect 835 4225 855 4245
rect 1075 4225 1095 4245
rect 1435 4225 1455 4245
rect 1675 4225 1695 4245
rect 1855 4225 1875 4245
rect 2035 4225 2055 4245
rect 2215 4225 2235 4245
rect 2395 4225 2415 4245
rect 2495 4225 2515 4245
rect 15 2720 35 2745
rect 115 2720 135 2745
rect 2395 2720 2415 2745
rect 2495 2720 2515 2745
rect 1185 1930 1210 1950
rect 1320 1930 1345 1950
rect 1280 1275 1300 1295
rect 15 1220 35 1245
rect 115 1220 135 1245
rect 295 1220 315 1245
rect 475 1220 495 1245
rect 655 1220 675 1245
rect 835 1220 855 1245
rect 1075 1220 1095 1245
rect 1435 1220 1455 1245
rect 1675 1220 1695 1245
rect 1855 1220 1875 1245
rect 2035 1220 2055 1245
rect 2215 1220 2235 1245
rect 2395 1220 2415 1245
rect 2495 1220 2515 1245
rect 1280 1115 1300 1135
<< locali >>
rect 1210 5820 2650 5840
rect 5 5745 45 5750
rect -35 5725 15 5745
rect 35 5725 45 5745
rect -35 5720 45 5725
rect 955 5745 995 5755
rect 955 5725 965 5745
rect 985 5725 995 5745
rect -35 5695 -15 5720
rect 955 5715 995 5725
rect 1065 5745 1105 5750
rect 1065 5725 1075 5745
rect 1095 5725 1145 5745
rect 1065 5720 1105 5725
rect -95 5685 -5 5695
rect -95 4515 -85 5685
rect -60 4515 -35 5685
rect -15 4515 -5 5685
rect -95 4505 -5 4515
rect 55 5685 95 5695
rect 55 4515 65 5685
rect 85 4515 95 5685
rect 55 4505 95 4515
rect 155 5685 195 5695
rect 155 4515 165 5685
rect 185 4515 195 5685
rect 155 4505 195 4515
rect 295 5685 335 5695
rect 295 4515 305 5685
rect 325 4515 335 5685
rect 295 4505 335 4515
rect 395 5685 435 5695
rect 395 4515 405 5685
rect 425 4515 435 5685
rect 395 4505 435 4515
rect 495 5685 535 5695
rect 495 4515 505 5685
rect 525 4515 535 5685
rect 495 4505 535 4515
rect 595 5685 635 5695
rect 595 4515 605 5685
rect 625 4515 635 5685
rect 595 4505 635 4515
rect 695 5685 735 5695
rect 695 4515 705 5685
rect 725 4525 735 5685
rect 725 4515 955 4525
rect 695 4505 955 4515
rect 175 4295 195 4505
rect 65 4275 805 4295
rect -25 4245 45 4250
rect -25 4225 15 4245
rect 35 4225 45 4245
rect -25 4215 45 4225
rect -25 4195 -5 4215
rect 65 4195 85 4275
rect 105 4245 145 4250
rect 105 4225 115 4245
rect 135 4225 185 4245
rect 105 4215 145 4225
rect 165 4195 185 4225
rect 245 4195 265 4275
rect 285 4245 325 4250
rect 285 4225 295 4245
rect 315 4225 365 4245
rect 285 4215 325 4225
rect 345 4195 365 4225
rect 425 4195 445 4275
rect 465 4245 505 4250
rect 465 4225 475 4245
rect 495 4225 545 4245
rect 465 4215 505 4225
rect 525 4195 545 4225
rect 605 4195 625 4275
rect 645 4245 685 4250
rect 645 4225 655 4245
rect 675 4225 725 4245
rect 645 4215 685 4225
rect 705 4195 725 4225
rect 785 4195 805 4275
rect 825 4245 905 4250
rect 825 4225 835 4245
rect 855 4225 905 4245
rect 825 4215 865 4225
rect 885 4195 905 4225
rect -95 4185 -5 4195
rect -95 3015 -85 4185
rect -60 3015 -35 4185
rect -15 3015 -5 4185
rect -95 3005 -5 3015
rect 55 4185 95 4195
rect 55 3015 65 4185
rect 85 3015 95 4185
rect 55 3005 95 3015
rect 155 4185 195 4195
rect 155 3015 165 4185
rect 185 3015 195 4185
rect 155 3005 195 3015
rect 235 4185 275 4195
rect 235 3015 245 4185
rect 265 3015 275 4185
rect 235 3005 275 3015
rect 335 4185 375 4195
rect 335 3015 345 4185
rect 365 3015 375 4185
rect 335 3005 375 3015
rect 415 4185 455 4195
rect 415 3015 425 4185
rect 445 3015 455 4185
rect 415 3005 455 3015
rect 515 4185 555 4195
rect 515 3015 525 4185
rect 545 3015 555 4185
rect 515 3005 555 3015
rect 595 4185 635 4195
rect 595 3015 605 4185
rect 625 3015 635 4185
rect 595 3005 635 3015
rect 695 4185 735 4195
rect 695 3015 705 4185
rect 725 3015 735 4185
rect 695 3005 735 3015
rect 775 4185 815 4195
rect 775 3015 785 4185
rect 805 3015 815 4185
rect 775 3005 815 3015
rect 875 4185 915 4195
rect 875 3015 885 4185
rect 905 3015 915 4185
rect 875 3005 915 3015
rect 165 2985 185 3005
rect 345 2985 365 3005
rect 525 2985 545 3005
rect 705 2985 725 3005
rect 165 2965 725 2985
rect -120 2770 90 2790
rect 70 2750 90 2770
rect -25 2745 45 2750
rect -25 2720 15 2745
rect 35 2720 45 2745
rect -25 2715 45 2720
rect 70 2745 145 2750
rect 70 2720 115 2745
rect 135 2720 145 2745
rect 70 2715 145 2720
rect -25 2695 -5 2715
rect 70 2695 90 2715
rect 305 2695 325 2965
rect 885 2695 905 3005
rect -95 2685 -5 2695
rect -95 1515 -85 2685
rect -60 1515 -35 2685
rect -15 1515 -5 2685
rect -95 1505 -5 1515
rect 55 2685 95 2695
rect 55 1515 65 2685
rect 85 1515 95 2685
rect 55 1505 95 1515
rect 155 2685 195 2695
rect 155 1515 165 2685
rect 185 1515 195 2685
rect 155 1505 195 1515
rect 295 2685 335 2695
rect 295 1515 305 2685
rect 325 1515 335 2685
rect 295 1505 335 1515
rect 395 2685 435 2695
rect 395 1515 405 2685
rect 425 1515 435 2685
rect 395 1505 435 1515
rect 495 2685 535 2695
rect 495 1515 505 2685
rect 525 1515 535 2685
rect 495 1505 535 1515
rect 595 2685 635 2695
rect 595 1515 605 2685
rect 625 1515 635 2685
rect 595 1505 635 1515
rect 695 2685 735 2695
rect 695 1515 705 2685
rect 725 1515 735 2685
rect 695 1505 735 1515
rect 775 2685 815 2695
rect 775 1515 785 2685
rect 805 1515 815 2685
rect 775 1505 815 1515
rect 875 2685 915 2695
rect 875 1515 885 2685
rect 905 1515 915 2685
rect 875 1505 915 1515
rect 935 1290 955 4505
rect 975 2825 995 5715
rect 1125 5695 1145 5725
rect 1015 5685 1055 5695
rect 1015 4515 1025 5685
rect 1045 4515 1055 5685
rect 1015 4505 1055 4515
rect 1115 5685 1155 5695
rect 1115 4515 1125 5685
rect 1145 4515 1155 5685
rect 1115 4505 1155 4515
rect 1065 4475 1105 4485
rect 1065 4455 1075 4475
rect 1095 4455 1105 4475
rect 1065 4450 1105 4455
rect 1075 4250 1095 4450
rect 1210 4345 1230 5820
rect 1290 5780 2650 5800
rect 1290 5770 1320 5780
rect 1280 5765 1320 5770
rect 1280 5745 1290 5765
rect 1310 5745 1320 5765
rect 1425 5745 1465 5750
rect 1280 5740 1320 5745
rect 1385 5725 1435 5745
rect 1455 5725 1465 5745
rect 1385 5695 1405 5725
rect 1425 5720 1465 5725
rect 1535 5745 1575 5755
rect 1535 5725 1545 5745
rect 1565 5725 1575 5745
rect 1535 5715 1575 5725
rect 2485 5745 2525 5750
rect 2485 5725 2495 5745
rect 2515 5725 2565 5745
rect 2485 5720 2565 5725
rect 1375 5685 1415 5695
rect 1375 4515 1385 5685
rect 1405 4515 1415 5685
rect 1375 4505 1415 4515
rect 1475 5685 1515 5695
rect 1475 4515 1485 5685
rect 1505 4515 1515 5685
rect 1475 4505 1515 4515
rect 1425 4475 1465 4485
rect 1425 4455 1435 4475
rect 1455 4455 1465 4475
rect 1425 4450 1465 4455
rect 1200 4340 1240 4345
rect 1200 4320 1210 4340
rect 1230 4320 1240 4340
rect 1200 4315 1240 4320
rect 1435 4250 1455 4450
rect 1065 4245 1105 4250
rect 1065 4225 1075 4245
rect 1095 4225 1105 4245
rect 1065 4215 1105 4225
rect 1425 4245 1465 4250
rect 1425 4225 1435 4245
rect 1455 4225 1465 4245
rect 1425 4215 1465 4225
rect 1015 4185 1055 4195
rect 1015 3015 1025 4185
rect 1045 3015 1055 4185
rect 1015 3005 1055 3015
rect 1115 4185 1155 4195
rect 1115 3015 1125 4185
rect 1145 3025 1155 4185
rect 1375 4185 1415 4195
rect 1375 3025 1385 4185
rect 1145 3015 1220 3025
rect 1115 3005 1220 3015
rect 975 2805 1045 2825
rect 1025 2695 1045 2805
rect 1015 2685 1055 2695
rect 1015 1515 1025 2685
rect 1045 1515 1055 2685
rect 1015 1505 1055 1515
rect 1115 2685 1155 2695
rect 1115 1515 1125 2685
rect 1145 1515 1155 2685
rect 1200 1955 1220 3005
rect 1175 1950 1220 1955
rect 1175 1930 1185 1950
rect 1210 1930 1220 1950
rect 1175 1925 1220 1930
rect 1310 3015 1385 3025
rect 1405 3015 1415 4185
rect 1310 3005 1415 3015
rect 1475 4185 1515 4195
rect 1475 3015 1485 4185
rect 1505 3015 1515 4185
rect 1475 3005 1515 3015
rect 1310 1955 1330 3005
rect 1535 2825 1555 5715
rect 2545 5695 2565 5720
rect 1795 5685 1835 5695
rect 1795 4525 1805 5685
rect 1485 2805 1555 2825
rect 1575 4515 1805 4525
rect 1825 4515 1835 5685
rect 1575 4505 1835 4515
rect 1895 5685 1935 5695
rect 1895 4515 1905 5685
rect 1925 4515 1935 5685
rect 1895 4505 1935 4515
rect 1995 5685 2035 5695
rect 1995 4515 2005 5685
rect 2025 4515 2035 5685
rect 1995 4505 2035 4515
rect 2095 5685 2135 5695
rect 2095 4515 2105 5685
rect 2125 4515 2135 5685
rect 2095 4505 2135 4515
rect 2195 5685 2235 5695
rect 2195 4515 2205 5685
rect 2225 4515 2235 5685
rect 2195 4505 2235 4515
rect 2335 5685 2375 5695
rect 2335 4515 2345 5685
rect 2365 4515 2375 5685
rect 2335 4505 2375 4515
rect 2435 5685 2475 5695
rect 2435 4515 2445 5685
rect 2465 4515 2475 5685
rect 2435 4505 2475 4515
rect 2535 5685 2625 5695
rect 2535 4515 2545 5685
rect 2565 4515 2590 5685
rect 2615 4515 2625 5685
rect 2535 4505 2625 4515
rect 1485 2695 1505 2805
rect 1375 2685 1415 2695
rect 1310 1950 1355 1955
rect 1310 1930 1320 1950
rect 1345 1930 1355 1950
rect 1310 1925 1355 1930
rect 1115 1505 1155 1515
rect 1375 1515 1385 2685
rect 1405 1515 1415 2685
rect 1375 1505 1415 1515
rect 1475 2685 1515 2695
rect 1475 1515 1485 2685
rect 1505 1515 1515 2685
rect 1475 1505 1515 1515
rect 1270 1295 1310 1305
rect 1270 1290 1280 1295
rect 935 1275 1280 1290
rect 1300 1290 1310 1295
rect 1575 1290 1595 4505
rect 2335 4295 2355 4505
rect 1725 4275 2465 4295
rect 1625 4245 1705 4250
rect 1625 4225 1675 4245
rect 1695 4225 1705 4245
rect 1625 4195 1645 4225
rect 1665 4215 1705 4225
rect 1725 4195 1745 4275
rect 1845 4245 1885 4250
rect 1805 4225 1855 4245
rect 1875 4225 1885 4245
rect 1805 4195 1825 4225
rect 1845 4215 1885 4225
rect 1905 4195 1925 4275
rect 2025 4245 2065 4250
rect 1985 4225 2035 4245
rect 2055 4225 2065 4245
rect 1985 4195 2005 4225
rect 2025 4215 2065 4225
rect 2085 4195 2105 4275
rect 2205 4245 2245 4250
rect 2165 4225 2215 4245
rect 2235 4225 2245 4245
rect 2165 4195 2185 4225
rect 2205 4215 2245 4225
rect 2265 4195 2285 4275
rect 2385 4245 2425 4250
rect 2345 4225 2395 4245
rect 2415 4225 2425 4245
rect 2345 4195 2365 4225
rect 2385 4215 2425 4225
rect 2445 4195 2465 4275
rect 2485 4245 2555 4250
rect 2485 4225 2495 4245
rect 2515 4225 2555 4245
rect 2485 4215 2555 4225
rect 2535 4195 2555 4215
rect 1615 4185 1655 4195
rect 1615 3015 1625 4185
rect 1645 3015 1655 4185
rect 1615 3005 1655 3015
rect 1715 4185 1755 4195
rect 1715 3015 1725 4185
rect 1745 3015 1755 4185
rect 1715 3005 1755 3015
rect 1795 4185 1835 4195
rect 1795 3015 1805 4185
rect 1825 3015 1835 4185
rect 1795 3005 1835 3015
rect 1895 4185 1935 4195
rect 1895 3015 1905 4185
rect 1925 3015 1935 4185
rect 1895 3005 1935 3015
rect 1975 4185 2015 4195
rect 1975 3015 1985 4185
rect 2005 3015 2015 4185
rect 1975 3005 2015 3015
rect 2075 4185 2115 4195
rect 2075 3015 2085 4185
rect 2105 3015 2115 4185
rect 2075 3005 2115 3015
rect 2155 4185 2195 4195
rect 2155 3015 2165 4185
rect 2185 3015 2195 4185
rect 2155 3005 2195 3015
rect 2255 4185 2295 4195
rect 2255 3015 2265 4185
rect 2285 3015 2295 4185
rect 2255 3005 2295 3015
rect 2335 4185 2375 4195
rect 2335 3015 2345 4185
rect 2365 3015 2375 4185
rect 2335 3005 2375 3015
rect 2435 4185 2475 4195
rect 2435 3015 2445 4185
rect 2465 3015 2475 4185
rect 2435 3005 2475 3015
rect 2535 4185 2625 4195
rect 2535 3015 2545 4185
rect 2565 3015 2590 4185
rect 2615 3015 2625 4185
rect 2535 3005 2625 3015
rect 1625 2695 1645 3005
rect 1805 2985 1825 3005
rect 1985 2985 2005 3005
rect 2165 2985 2185 3005
rect 2345 2985 2365 3005
rect 1805 2965 2365 2985
rect 2205 2695 2225 2965
rect 2385 2745 2460 2750
rect 2385 2720 2395 2745
rect 2415 2720 2460 2745
rect 2385 2715 2460 2720
rect 2485 2745 2555 2750
rect 2485 2720 2495 2745
rect 2515 2720 2555 2745
rect 2485 2715 2555 2720
rect 2440 2695 2460 2715
rect 2535 2695 2555 2715
rect 1615 2685 1655 2695
rect 1615 1515 1625 2685
rect 1645 1515 1655 2685
rect 1615 1505 1655 1515
rect 1715 2685 1755 2695
rect 1715 1515 1725 2685
rect 1745 1515 1755 2685
rect 1715 1505 1755 1515
rect 1795 2685 1835 2695
rect 1795 1515 1805 2685
rect 1825 1515 1835 2685
rect 1795 1505 1835 1515
rect 1895 2685 1935 2695
rect 1895 1515 1905 2685
rect 1925 1515 1935 2685
rect 1895 1505 1935 1515
rect 1995 2685 2035 2695
rect 1995 1515 2005 2685
rect 2025 1515 2035 2685
rect 1995 1505 2035 1515
rect 2095 2685 2135 2695
rect 2095 1515 2105 2685
rect 2125 1515 2135 2685
rect 2095 1505 2135 1515
rect 2195 2685 2235 2695
rect 2195 1515 2205 2685
rect 2225 1515 2235 2685
rect 2195 1505 2235 1515
rect 2335 2685 2375 2695
rect 2335 1515 2345 2685
rect 2365 1515 2375 2685
rect 2335 1505 2375 1515
rect 2435 2685 2475 2695
rect 2435 1515 2445 2685
rect 2465 1515 2475 2685
rect 2435 1505 2475 1515
rect 2535 2685 2625 2695
rect 2535 1515 2545 2685
rect 2565 1515 2590 2685
rect 2615 1515 2625 2685
rect 2535 1505 2625 1515
rect 1300 1275 1595 1290
rect 935 1270 1595 1275
rect 935 1250 955 1270
rect 1270 1265 1310 1270
rect 1575 1250 1595 1270
rect 5 1245 45 1250
rect -35 1220 15 1245
rect 35 1220 45 1245
rect -35 1195 -15 1220
rect 5 1215 45 1220
rect 105 1245 145 1250
rect 285 1245 325 1250
rect 465 1245 505 1250
rect 645 1245 685 1250
rect 825 1245 955 1250
rect 105 1220 115 1245
rect 135 1220 185 1245
rect 105 1215 145 1220
rect 165 1195 185 1220
rect 285 1220 295 1245
rect 315 1220 365 1245
rect 285 1215 325 1220
rect 345 1195 365 1220
rect 465 1220 475 1245
rect 495 1220 545 1245
rect 465 1215 505 1220
rect 525 1195 545 1220
rect 645 1220 655 1245
rect 675 1220 725 1245
rect 645 1215 685 1220
rect 705 1195 725 1220
rect 825 1220 835 1245
rect 855 1230 955 1245
rect 1065 1245 1105 1250
rect 855 1220 865 1230
rect 825 1215 865 1220
rect 1065 1220 1075 1245
rect 1095 1240 1105 1245
rect 1425 1245 1465 1250
rect 1425 1240 1435 1245
rect 1095 1220 1435 1240
rect 1455 1220 1465 1245
rect 1575 1245 1705 1250
rect 1845 1245 1885 1250
rect 2025 1245 2065 1250
rect 2205 1245 2245 1250
rect 2385 1245 2425 1250
rect 1575 1230 1675 1245
rect 1065 1215 1105 1220
rect 1125 1195 1145 1220
rect -95 1185 -5 1195
rect -95 15 -85 1185
rect -60 15 -35 1185
rect -15 15 -5 1185
rect -95 5 -5 15
rect 55 1185 95 1195
rect 55 15 65 1185
rect 85 15 95 1185
rect 55 5 95 15
rect 155 1185 195 1195
rect 155 15 165 1185
rect 185 15 195 1185
rect 155 5 195 15
rect 235 1185 275 1195
rect 235 15 245 1185
rect 265 15 275 1185
rect 235 5 275 15
rect 335 1185 375 1195
rect 335 15 345 1185
rect 365 15 375 1185
rect 335 5 375 15
rect 415 1185 455 1195
rect 415 15 425 1185
rect 445 15 455 1185
rect 415 5 455 15
rect 515 1185 555 1195
rect 515 15 525 1185
rect 545 15 555 1185
rect 515 5 555 15
rect 595 1185 635 1195
rect 595 15 605 1185
rect 625 15 635 1185
rect 595 5 635 15
rect 695 1185 735 1195
rect 695 15 705 1185
rect 725 15 735 1185
rect 695 5 735 15
rect 775 1185 815 1195
rect 775 15 785 1185
rect 805 15 815 1185
rect 775 5 815 15
rect 875 1185 915 1195
rect 875 15 885 1185
rect 905 15 915 1185
rect 875 5 915 15
rect 1015 1185 1055 1195
rect 1015 15 1025 1185
rect 1045 15 1055 1185
rect 1015 5 1055 15
rect 1115 1185 1155 1195
rect 1115 15 1125 1185
rect 1145 15 1155 1185
rect 1115 5 1155 15
rect 75 -15 95 5
rect 235 -15 255 5
rect 415 -15 435 5
rect 595 -15 615 5
rect 875 -15 895 5
rect 1015 -15 1035 5
rect 75 -35 1035 -15
rect 1225 -100 1245 1220
rect 1385 1195 1405 1220
rect 1425 1215 1465 1220
rect 1665 1220 1675 1230
rect 1695 1220 1705 1245
rect 1665 1215 1705 1220
rect 1805 1220 1855 1245
rect 1875 1220 1885 1245
rect 1805 1195 1825 1220
rect 1845 1215 1885 1220
rect 1985 1220 2035 1245
rect 2055 1220 2065 1245
rect 1985 1195 2005 1220
rect 2025 1215 2065 1220
rect 2165 1220 2215 1245
rect 2235 1220 2245 1245
rect 2165 1195 2185 1220
rect 2205 1215 2245 1220
rect 2345 1220 2395 1245
rect 2415 1220 2425 1245
rect 2345 1195 2365 1220
rect 2385 1215 2425 1220
rect 2485 1245 2525 1250
rect 2485 1220 2495 1245
rect 2515 1220 2565 1245
rect 2485 1215 2525 1220
rect 2545 1195 2565 1220
rect 1375 1185 1415 1195
rect 1270 1135 1310 1145
rect 1270 1115 1280 1135
rect 1300 1115 1310 1135
rect 1270 1105 1310 1115
rect 1275 -55 1295 1105
rect 1375 15 1385 1185
rect 1405 15 1415 1185
rect 1375 5 1415 15
rect 1475 1185 1515 1195
rect 1475 15 1485 1185
rect 1505 15 1515 1185
rect 1475 5 1515 15
rect 1615 1185 1655 1195
rect 1615 15 1625 1185
rect 1645 15 1655 1185
rect 1615 5 1655 15
rect 1715 1185 1755 1195
rect 1715 15 1725 1185
rect 1745 15 1755 1185
rect 1715 5 1755 15
rect 1795 1185 1835 1195
rect 1795 15 1805 1185
rect 1825 15 1835 1185
rect 1795 5 1835 15
rect 1895 1185 1935 1195
rect 1895 15 1905 1185
rect 1925 15 1935 1185
rect 1895 5 1935 15
rect 1975 1185 2015 1195
rect 1975 15 1985 1185
rect 2005 15 2015 1185
rect 1975 5 2015 15
rect 2075 1185 2115 1195
rect 2075 15 2085 1185
rect 2105 15 2115 1185
rect 2075 5 2115 15
rect 2155 1185 2195 1195
rect 2155 15 2165 1185
rect 2185 15 2195 1185
rect 2155 5 2195 15
rect 2255 1185 2295 1195
rect 2255 15 2265 1185
rect 2285 15 2295 1185
rect 2255 5 2295 15
rect 2335 1185 2375 1195
rect 2335 15 2345 1185
rect 2365 15 2375 1185
rect 2335 5 2375 15
rect 2435 1185 2475 1195
rect 2435 15 2445 1185
rect 2465 15 2475 1185
rect 2435 5 2475 15
rect 2535 1185 2625 1195
rect 2535 15 2545 1185
rect 2565 15 2590 1185
rect 2615 15 2625 1185
rect 2535 5 2625 15
rect 1495 -15 1515 5
rect 1635 -15 1655 5
rect 1915 -15 1935 5
rect 2095 -15 2115 5
rect 2275 -15 2295 5
rect 2435 -15 2455 5
rect 1495 -35 2455 -15
rect 1275 -75 2650 -55
rect 1225 -120 2650 -100
<< viali >>
rect -85 4515 -60 5685
rect -35 4515 -15 5685
rect 65 4515 85 5685
rect 305 4515 325 5685
rect -85 3015 -60 4185
rect -35 3015 -15 4185
rect -85 1515 -60 2685
rect -35 1515 -15 2685
rect 165 1515 185 2685
rect 705 1515 725 2685
rect 785 1515 805 2685
rect 1025 4515 1045 5685
rect 1485 4515 1505 5685
rect 1025 3015 1045 4185
rect 1125 1515 1145 2685
rect 1485 3015 1505 4185
rect 2205 4515 2225 5685
rect 2445 4515 2465 5685
rect 2545 4515 2565 5685
rect 2590 4515 2615 5685
rect 1385 1515 1405 2685
rect 2545 3015 2565 4185
rect 2590 3015 2615 4185
rect 1725 1515 1745 2685
rect 1805 1515 1825 2685
rect 2345 1515 2365 2685
rect 2545 1515 2565 2685
rect 2590 1515 2615 2685
rect -85 15 -60 1185
rect -35 15 -15 1185
rect 785 15 805 1185
rect 1725 15 1745 1185
rect 2545 15 2565 1185
rect 2590 15 2615 1185
<< metal1 >>
rect -120 5685 2650 5700
rect -120 4515 -85 5685
rect -60 4515 -35 5685
rect -15 4515 65 5685
rect 85 4515 305 5685
rect 325 4515 1025 5685
rect 1045 4515 1485 5685
rect 1505 4515 2205 5685
rect 2225 4515 2445 5685
rect 2465 4515 2545 5685
rect 2565 4515 2590 5685
rect 2615 4515 2650 5685
rect -120 4185 2650 4515
rect -120 3015 -85 4185
rect -60 3015 -35 4185
rect -15 3015 1025 4185
rect 1045 3015 1485 4185
rect 1505 3015 2545 4185
rect 2565 3015 2590 4185
rect 2615 3015 2650 4185
rect -120 3000 2650 3015
rect -120 2685 2650 2700
rect -120 1515 -85 2685
rect -60 1515 -35 2685
rect -15 1515 165 2685
rect 185 1515 705 2685
rect 725 1515 785 2685
rect 805 1515 1125 2685
rect 1145 1515 1385 2685
rect 1405 1515 1725 2685
rect 1745 1515 1805 2685
rect 1825 1515 2345 2685
rect 2365 1515 2545 2685
rect 2565 1515 2590 2685
rect 2615 1515 2650 2685
rect -120 1185 2650 1515
rect -120 15 -85 1185
rect -60 15 -35 1185
rect -15 15 785 1185
rect 805 15 1725 1185
rect 1745 15 2545 1185
rect 2565 15 2590 1185
rect 2615 15 2650 1185
rect -120 5 2650 15
rect -100 0 2650 5
<< labels >>
rlabel locali -120 2780 -120 2780 7 VB
port 1 w
rlabel metal1 -120 3015 -120 3015 7 VP
port 2 w
rlabel metal1 -120 2685 -120 2685 7 VN
port 3 w
rlabel locali 2650 5830 2650 5830 3 VCP
port 4 e
rlabel locali 2650 5790 2650 5790 3 VBP
port 5 e
rlabel locali 2650 -65 2650 -65 3 VBN
port 6 e
rlabel locali 2650 -110 2650 -110 3 VCN
port 7 e
<< end >>
