magic
tech sky130A
timestamp 1695854801
<< nwell >>
rect -35 1195 195 2280
<< nmos >>
rect 105 1010 120 1110
<< pmos >>
rect 105 1345 120 1445
<< ndiff >>
rect 55 1095 105 1110
rect 55 1025 70 1095
rect 90 1025 105 1095
rect 55 1010 105 1025
rect 120 1095 170 1110
rect 120 1025 135 1095
rect 155 1025 170 1095
rect 120 1010 170 1025
<< pdiff >>
rect 55 1430 105 1445
rect 55 1360 70 1430
rect 90 1360 105 1430
rect 55 1345 105 1360
rect 120 1430 170 1445
rect 120 1360 135 1430
rect 155 1360 170 1430
rect 120 1345 170 1360
<< ndiffc >>
rect 70 1025 90 1095
rect 135 1025 155 1095
<< pdiffc >>
rect 70 1360 90 1430
rect 135 1360 155 1430
<< psubdiff >>
rect 5 1095 55 1110
rect 5 1025 20 1095
rect 40 1025 55 1095
rect 5 1010 55 1025
<< nsubdiff >>
rect 5 1430 55 1445
rect 5 1360 20 1430
rect 40 1360 55 1430
rect 5 1345 55 1360
<< psubdiffcont >>
rect 20 1025 40 1095
<< nsubdiffcont >>
rect 20 1360 40 1430
<< poly >>
rect 105 1445 120 1460
rect 105 1110 120 1345
rect 105 995 120 1010
rect 105 985 145 995
rect 105 965 115 985
rect 135 965 145 985
rect 105 955 145 965
<< polycont >>
rect 115 965 135 985
<< locali >>
rect 10 1430 100 1440
rect 10 1360 20 1430
rect 40 1360 70 1430
rect 90 1360 100 1430
rect 10 1350 100 1360
rect 125 1430 165 1440
rect 125 1360 135 1430
rect 155 1360 165 1430
rect 125 1350 165 1360
rect 145 1325 165 1350
rect 145 1295 195 1325
rect 145 1105 165 1295
rect 10 1095 100 1105
rect 10 1025 20 1095
rect 40 1025 70 1095
rect 90 1025 100 1095
rect 10 1015 100 1025
rect 125 1095 165 1105
rect 125 1025 135 1095
rect 155 1025 165 1095
rect 125 1015 165 1025
rect -35 985 145 995
rect -35 965 115 985
rect 135 965 145 985
rect 105 955 145 965
<< viali >>
rect 20 1360 40 1430
rect 70 1360 90 1430
rect 20 1025 40 1095
rect 70 1025 90 1095
<< metal1 >>
rect -35 1430 195 2265
rect -35 1360 20 1430
rect 40 1360 70 1430
rect 90 1360 195 1430
rect -35 1225 195 1360
rect -35 1095 195 1120
rect -35 1025 20 1095
rect 40 1025 70 1095
rect 90 1025 195 1095
rect -35 90 195 1025
<< labels >>
rlabel metal1 -35 1610 -35 1610 7 VP
port 3 w
rlabel metal1 -35 865 -35 865 7 VN
port 4 w
rlabel locali 195 1310 195 1310 3 Y
port 2 e
rlabel locali -35 980 -35 980 7 A
port 1 w
<< end >>
